----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 07.11.2022 19:01:24
-- Design Name: 
-- Module Name: layer_template - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity layer is
    Port ( 
        x : in STD_LOGIC_VECTOR;
        y : out STD_LOGIC_VECTOR
   );
end layer;

architecture layer_1 of layer is

    Component perceptron
    Generic (
        WEIGHTS : STD_LOGIC_VECTOR := (others => '0');
        SHIFT : Integer;     -- number of shift (left + or right -)
        B : Integer;          -- bias of batch norm
        BATCH_POSITIVE : Boolean    
    );
    Port ( 
        x : in STD_LOGIC_VECTOR;
        y : out STD_LOGIC_VECTOR
   );
    end component;
    
    -- Signals
    signal p0_in : STD_LOGIC_VECTOR(0 to 36 - 1);
	signal p0_out : STD_LOGIC;
	signal p1_in : STD_LOGIC_VECTOR(0 to 117 - 1);
	signal p1_out : STD_LOGIC;
	signal p2_in : STD_LOGIC_VECTOR(0 to 138 - 1);
	signal p2_out : STD_LOGIC;
	signal p3_in : STD_LOGIC_VECTOR(0 to 71 - 1);
	signal p3_out : STD_LOGIC;
	signal p4_in : STD_LOGIC_VECTOR(0 to 89 - 1);
	signal p4_out : STD_LOGIC;
	signal p5_in : STD_LOGIC_VECTOR(0 to 47 - 1);
	signal p5_out : STD_LOGIC;
	signal p6_in : STD_LOGIC_VECTOR(0 to 104 - 1);
	signal p6_out : STD_LOGIC;
	signal p7_in : STD_LOGIC_VECTOR(0 to 85 - 1);
	signal p7_out : STD_LOGIC;
	signal p8_in : STD_LOGIC_VECTOR(0 to 42 - 1);
	signal p8_out : STD_LOGIC;
	signal p9_in : STD_LOGIC_VECTOR(0 to 75 - 1);
	signal p9_out : STD_LOGIC;
	signal p10_in : STD_LOGIC_VECTOR(0 to 96 - 1);
	signal p10_out : STD_LOGIC;
	signal p11_in : STD_LOGIC_VECTOR(0 to 103 - 1);
	signal p11_out : STD_LOGIC;
	signal p12_in : STD_LOGIC_VECTOR(0 to 94 - 1);
	signal p12_out : STD_LOGIC;
	signal p13_in : STD_LOGIC_VECTOR(0 to 59 - 1);
	signal p13_out : STD_LOGIC;
	signal p14_in : STD_LOGIC_VECTOR(0 to 117 - 1);
	signal p14_out : STD_LOGIC;
	signal p15_in : STD_LOGIC_VECTOR(0 to 104 - 1);
	signal p15_out : STD_LOGIC;
	signal p16_in : STD_LOGIC_VECTOR(0 to 84 - 1);
	signal p16_out : STD_LOGIC;
	signal p17_in : STD_LOGIC_VECTOR(0 to 68 - 1);
	signal p17_out : STD_LOGIC;
	signal p18_in : STD_LOGIC_VECTOR(0 to 121 - 1);
	signal p18_out : STD_LOGIC;
	signal p19_in : STD_LOGIC_VECTOR(0 to 92 - 1);
	signal p19_out : STD_LOGIC;
	signal p20_in : STD_LOGIC_VECTOR(0 to 121 - 1);
	signal p20_out : STD_LOGIC;
	signal p21_in : STD_LOGIC_VECTOR(0 to 63 - 1);
	signal p21_out : STD_LOGIC;
	signal p22_in : STD_LOGIC_VECTOR(0 to 80 - 1);
	signal p22_out : STD_LOGIC;
	signal p23_in : STD_LOGIC_VECTOR(0 to 135 - 1);
	signal p23_out : STD_LOGIC;
	signal p24_in : STD_LOGIC_VECTOR(0 to 53 - 1);
	signal p24_out : STD_LOGIC;
	signal p25_in : STD_LOGIC_VECTOR(0 to 93 - 1);
	signal p25_out : STD_LOGIC;
	signal p26_in : STD_LOGIC_VECTOR(0 to 76 - 1);
	signal p26_out : STD_LOGIC;
	signal p27_in : STD_LOGIC_VECTOR(0 to 94 - 1);
	signal p27_out : STD_LOGIC;
	signal p28_in : STD_LOGIC_VECTOR(0 to 103 - 1);
	signal p28_out : STD_LOGIC;
	signal p29_in : STD_LOGIC_VECTOR(0 to 64 - 1);
	signal p29_out : STD_LOGIC;
	signal p30_in : STD_LOGIC_VECTOR(0 to 121 - 1);
	signal p30_out : STD_LOGIC;
	signal p31_in : STD_LOGIC_VECTOR(0 to 96 - 1);
	signal p31_out : STD_LOGIC;
	signal p32_in : STD_LOGIC_VECTOR(0 to 80 - 1);
	signal p32_out : STD_LOGIC;
	signal p33_in : STD_LOGIC_VECTOR(0 to 213 - 1);
	signal p33_out : STD_LOGIC;
	signal p34_in : STD_LOGIC_VECTOR(0 to 149 - 1);
	signal p34_out : STD_LOGIC;
	signal p35_in : STD_LOGIC_VECTOR(0 to 209 - 1);
	signal p35_out : STD_LOGIC;
	signal p36_in : STD_LOGIC_VECTOR(0 to 116 - 1);
	signal p36_out : STD_LOGIC;
	signal p37_in : STD_LOGIC_VECTOR(0 to 114 - 1);
	signal p37_out : STD_LOGIC;
	signal p38_in : STD_LOGIC_VECTOR(0 to 75 - 1);
	signal p38_out : STD_LOGIC;
	signal p39_in : STD_LOGIC_VECTOR(0 to 100 - 1);
	signal p39_out : STD_LOGIC;
	signal p40_in : STD_LOGIC_VECTOR(0 to 89 - 1);
	signal p40_out : STD_LOGIC;
	signal p41_in : STD_LOGIC_VECTOR(0 to 87 - 1);
	signal p41_out : STD_LOGIC;
	signal p42_in : STD_LOGIC_VECTOR(0 to 122 - 1);
	signal p42_out : STD_LOGIC;
	signal p43_in : STD_LOGIC_VECTOR(0 to 101 - 1);
	signal p43_out : STD_LOGIC;
	signal p44_in : STD_LOGIC_VECTOR(0 to 98 - 1);
	signal p44_out : STD_LOGIC;
	signal p45_in : STD_LOGIC_VECTOR(0 to 104 - 1);
	signal p45_out : STD_LOGIC;
	signal p46_in : STD_LOGIC_VECTOR(0 to 124 - 1);
	signal p46_out : STD_LOGIC;
	signal p47_in : STD_LOGIC_VECTOR(0 to 64 - 1);
	signal p47_out : STD_LOGIC;
	signal p48_in : STD_LOGIC_VECTOR(0 to 120 - 1);
	signal p48_out : STD_LOGIC;
	signal p49_in : STD_LOGIC_VECTOR(0 to 88 - 1);
	signal p49_out : STD_LOGIC;
	signal p50_in : STD_LOGIC_VECTOR(0 to 94 - 1);
	signal p50_out : STD_LOGIC;
	signal p51_in : STD_LOGIC_VECTOR(0 to 104 - 1);
	signal p51_out : STD_LOGIC;
	signal p52_in : STD_LOGIC_VECTOR(0 to 85 - 1);
	signal p52_out : STD_LOGIC;
	signal p53_in : STD_LOGIC_VECTOR(0 to 80 - 1);
	signal p53_out : STD_LOGIC;
	signal p54_in : STD_LOGIC_VECTOR(0 to 85 - 1);
	signal p54_out : STD_LOGIC;
	signal p55_in : STD_LOGIC_VECTOR(0 to 67 - 1);
	signal p55_out : STD_LOGIC;
	signal p56_in : STD_LOGIC_VECTOR(0 to 107 - 1);
	signal p56_out : STD_LOGIC;
	signal p57_in : STD_LOGIC_VECTOR(0 to 79 - 1);
	signal p57_out : STD_LOGIC;
	signal p58_in : STD_LOGIC_VECTOR(0 to 64 - 1);
	signal p58_out : STD_LOGIC;
	signal p59_in : STD_LOGIC_VECTOR(0 to 109 - 1);
	signal p59_out : STD_LOGIC;
	signal p60_in : STD_LOGIC_VECTOR(0 to 129 - 1);
	signal p60_out : STD_LOGIC;
	signal p61_in : STD_LOGIC_VECTOR(0 to 136 - 1);
	signal p61_out : STD_LOGIC;
	signal p62_in : STD_LOGIC_VECTOR(0 to 73 - 1);
	signal p62_out : STD_LOGIC;
	signal p63_in : STD_LOGIC_VECTOR(0 to 193 - 1);
	signal p63_out : STD_LOGIC;
	signal p64_in : STD_LOGIC_VECTOR(0 to 159 - 1);
	signal p64_out : STD_LOGIC;
	signal p65_in : STD_LOGIC_VECTOR(0 to 66 - 1);
	signal p65_out : STD_LOGIC;
	signal p66_in : STD_LOGIC_VECTOR(0 to 110 - 1);
	signal p66_out : STD_LOGIC;
	signal p67_in : STD_LOGIC_VECTOR(0 to 51 - 1);
	signal p67_out : STD_LOGIC;
	signal p68_in : STD_LOGIC_VECTOR(0 to 68 - 1);
	signal p68_out : STD_LOGIC;
	signal p69_in : STD_LOGIC_VECTOR(0 to 76 - 1);
	signal p69_out : STD_LOGIC;
	signal p70_in : STD_LOGIC_VECTOR(0 to 86 - 1);
	signal p70_out : STD_LOGIC;
	signal p71_in : STD_LOGIC_VECTOR(0 to 96 - 1);
	signal p71_out : STD_LOGIC;
	signal p72_in : STD_LOGIC_VECTOR(0 to 68 - 1);
	signal p72_out : STD_LOGIC;
	signal p73_in : STD_LOGIC_VECTOR(0 to 45 - 1);
	signal p73_out : STD_LOGIC;
	signal p74_in : STD_LOGIC_VECTOR(0 to 78 - 1);
	signal p74_out : STD_LOGIC;
	signal p75_in : STD_LOGIC_VECTOR(0 to 86 - 1);
	signal p75_out : STD_LOGIC;
	signal p76_in : STD_LOGIC_VECTOR(0 to 78 - 1);
	signal p76_out : STD_LOGIC;
	signal p77_in : STD_LOGIC_VECTOR(0 to 91 - 1);
	signal p77_out : STD_LOGIC;
	signal p78_in : STD_LOGIC_VECTOR(0 to 73 - 1);
	signal p78_out : STD_LOGIC;
	signal p79_in : STD_LOGIC_VECTOR(0 to 69 - 1);
	signal p79_out : STD_LOGIC;
	signal p80_in : STD_LOGIC_VECTOR(0 to 66 - 1);
	signal p80_out : STD_LOGIC;
	signal p81_in : STD_LOGIC_VECTOR(0 to 99 - 1);
	signal p81_out : STD_LOGIC;
	signal p82_in : STD_LOGIC_VECTOR(0 to 98 - 1);
	signal p82_out : STD_LOGIC;
	signal p83_in : STD_LOGIC_VECTOR(0 to 106 - 1);
	signal p83_out : STD_LOGIC;
	signal p84_in : STD_LOGIC_VECTOR(0 to 130 - 1);
	signal p84_out : STD_LOGIC;
	signal p85_in : STD_LOGIC_VECTOR(0 to 93 - 1);
	signal p85_out : STD_LOGIC;
	signal p86_in : STD_LOGIC_VECTOR(0 to 85 - 1);
	signal p86_out : STD_LOGIC;
	signal p87_in : STD_LOGIC_VECTOR(0 to 106 - 1);
	signal p87_out : STD_LOGIC;
	signal p88_in : STD_LOGIC_VECTOR(0 to 72 - 1);
	signal p88_out : STD_LOGIC;
	signal p89_in : STD_LOGIC_VECTOR(0 to 129 - 1);
	signal p89_out : STD_LOGIC;
	signal p90_in : STD_LOGIC_VECTOR(0 to 84 - 1);
	signal p90_out : STD_LOGIC;
	signal p91_in : STD_LOGIC_VECTOR(0 to 118 - 1);
	signal p91_out : STD_LOGIC;
	signal p92_in : STD_LOGIC_VECTOR(0 to 87 - 1);
	signal p92_out : STD_LOGIC;
	signal p93_in : STD_LOGIC_VECTOR(0 to 93 - 1);
	signal p93_out : STD_LOGIC;
	signal p94_in : STD_LOGIC_VECTOR(0 to 80 - 1);
	signal p94_out : STD_LOGIC;
	signal p95_in : STD_LOGIC_VECTOR(0 to 80 - 1);
	signal p95_out : STD_LOGIC;
	signal p96_in : STD_LOGIC_VECTOR(0 to 135 - 1);
	signal p96_out : STD_LOGIC;
	signal p97_in : STD_LOGIC_VECTOR(0 to 159 - 1);
	signal p97_out : STD_LOGIC;
	signal p98_in : STD_LOGIC_VECTOR(0 to 119 - 1);
	signal p98_out : STD_LOGIC;
	signal p99_in : STD_LOGIC_VECTOR(0 to 121 - 1);
	signal p99_out : STD_LOGIC;
	signal p100_in : STD_LOGIC_VECTOR(0 to 94 - 1);
	signal p100_out : STD_LOGIC;
	signal p101_in : STD_LOGIC_VECTOR(0 to 100 - 1);
	signal p101_out : STD_LOGIC;
	signal p102_in : STD_LOGIC_VECTOR(0 to 81 - 1);
	signal p102_out : STD_LOGIC;
	signal p103_in : STD_LOGIC_VECTOR(0 to 122 - 1);
	signal p103_out : STD_LOGIC;
	signal p104_in : STD_LOGIC_VECTOR(0 to 126 - 1);
	signal p104_out : STD_LOGIC;
	signal p105_in : STD_LOGIC_VECTOR(0 to 84 - 1);
	signal p105_out : STD_LOGIC;
	signal p106_in : STD_LOGIC_VECTOR(0 to 78 - 1);
	signal p106_out : STD_LOGIC;
	signal p107_in : STD_LOGIC_VECTOR(0 to 178 - 1);
	signal p107_out : STD_LOGIC;
	signal p108_in : STD_LOGIC_VECTOR(0 to 70 - 1);
	signal p108_out : STD_LOGIC;
	signal p109_in : STD_LOGIC_VECTOR(0 to 58 - 1);
	signal p109_out : STD_LOGIC;
	signal p110_in : STD_LOGIC_VECTOR(0 to 107 - 1);
	signal p110_out : STD_LOGIC;
	signal p111_in : STD_LOGIC_VECTOR(0 to 134 - 1);
	signal p111_out : STD_LOGIC;
	signal p112_in : STD_LOGIC_VECTOR(0 to 83 - 1);
	signal p112_out : STD_LOGIC;
	signal p113_in : STD_LOGIC_VECTOR(0 to 95 - 1);
	signal p113_out : STD_LOGIC;
	signal p114_in : STD_LOGIC_VECTOR(0 to 77 - 1);
	signal p114_out : STD_LOGIC;
	signal p115_in : STD_LOGIC_VECTOR(0 to 69 - 1);
	signal p115_out : STD_LOGIC;
	signal p116_in : STD_LOGIC_VECTOR(0 to 122 - 1);
	signal p116_out : STD_LOGIC;
	signal p117_in : STD_LOGIC_VECTOR(0 to 181 - 1);
	signal p117_out : STD_LOGIC;
	signal p118_in : STD_LOGIC_VECTOR(0 to 196 - 1);
	signal p118_out : STD_LOGIC;
	signal p119_in : STD_LOGIC_VECTOR(0 to 105 - 1);
	signal p119_out : STD_LOGIC;
	signal p120_in : STD_LOGIC_VECTOR(0 to 49 - 1);
	signal p120_out : STD_LOGIC;
	signal p121_in : STD_LOGIC_VECTOR(0 to 99 - 1);
	signal p121_out : STD_LOGIC;
	signal p122_in : STD_LOGIC_VECTOR(0 to 134 - 1);
	signal p122_out : STD_LOGIC;
	signal p123_in : STD_LOGIC_VECTOR(0 to 105 - 1);
	signal p123_out : STD_LOGIC;
	signal p124_in : STD_LOGIC_VECTOR(0 to 55 - 1);
	signal p124_out : STD_LOGIC;
	signal p125_in : STD_LOGIC_VECTOR(0 to 120 - 1);
	signal p125_out : STD_LOGIC;
	signal p126_in : STD_LOGIC_VECTOR(0 to 135 - 1);
	signal p126_out : STD_LOGIC;
	signal p127_in : STD_LOGIC_VECTOR(0 to 67 - 1);
	signal p127_out : STD_LOGIC;
	signal p128_in : STD_LOGIC_VECTOR(0 to 81 - 1);
	signal p128_out : STD_LOGIC;
	signal p129_in : STD_LOGIC_VECTOR(0 to 100 - 1);
	signal p129_out : STD_LOGIC;
	signal p130_in : STD_LOGIC_VECTOR(0 to 94 - 1);
	signal p130_out : STD_LOGIC;
	signal p131_in : STD_LOGIC_VECTOR(0 to 60 - 1);
	signal p131_out : STD_LOGIC;
	signal p132_in : STD_LOGIC_VECTOR(0 to 79 - 1);
	signal p132_out : STD_LOGIC;
	signal p133_in : STD_LOGIC_VECTOR(0 to 99 - 1);
	signal p133_out : STD_LOGIC;
	signal p134_in : STD_LOGIC_VECTOR(0 to 121 - 1);
	signal p134_out : STD_LOGIC;
	signal p135_in : STD_LOGIC_VECTOR(0 to 98 - 1);
	signal p135_out : STD_LOGIC;
	signal p136_in : STD_LOGIC_VECTOR(0 to 72 - 1);
	signal p136_out : STD_LOGIC;
	signal p137_in : STD_LOGIC_VECTOR(0 to 70 - 1);
	signal p137_out : STD_LOGIC;
	signal p138_in : STD_LOGIC_VECTOR(0 to 116 - 1);
	signal p138_out : STD_LOGIC;
	signal p139_in : STD_LOGIC_VECTOR(0 to 98 - 1);
	signal p139_out : STD_LOGIC;
	signal p140_in : STD_LOGIC_VECTOR(0 to 82 - 1);
	signal p140_out : STD_LOGIC;
	signal p141_in : STD_LOGIC_VECTOR(0 to 76 - 1);
	signal p141_out : STD_LOGIC;
	signal p142_in : STD_LOGIC_VECTOR(0 to 182 - 1);
	signal p142_out : STD_LOGIC;
	signal p143_in : STD_LOGIC_VECTOR(0 to 72 - 1);
	signal p143_out : STD_LOGIC;
	signal p144_in : STD_LOGIC_VECTOR(0 to 114 - 1);
	signal p144_out : STD_LOGIC;
	signal p145_in : STD_LOGIC_VECTOR(0 to 92 - 1);
	signal p145_out : STD_LOGIC;
	signal p146_in : STD_LOGIC_VECTOR(0 to 82 - 1);
	signal p146_out : STD_LOGIC;
	signal p147_in : STD_LOGIC_VECTOR(0 to 237 - 1);
	signal p147_out : STD_LOGIC;
	signal p148_in : STD_LOGIC_VECTOR(0 to 118 - 1);
	signal p148_out : STD_LOGIC;
	signal p149_in : STD_LOGIC_VECTOR(0 to 188 - 1);
	signal p149_out : STD_LOGIC;
	signal p150_in : STD_LOGIC_VECTOR(0 to 142 - 1);
	signal p150_out : STD_LOGIC;
	signal p151_in : STD_LOGIC_VECTOR(0 to 120 - 1);
	signal p151_out : STD_LOGIC;
	signal p152_in : STD_LOGIC_VECTOR(0 to 137 - 1);
	signal p152_out : STD_LOGIC;
	signal p153_in : STD_LOGIC_VECTOR(0 to 43 - 1);
	signal p153_out : STD_LOGIC;
	signal p154_in : STD_LOGIC_VECTOR(0 to 172 - 1);
	signal p154_out : STD_LOGIC;
	signal p155_in : STD_LOGIC_VECTOR(0 to 117 - 1);
	signal p155_out : STD_LOGIC;
	signal p156_in : STD_LOGIC_VECTOR(0 to 116 - 1);
	signal p156_out : STD_LOGIC;
	signal p157_in : STD_LOGIC_VECTOR(0 to 145 - 1);
	signal p157_out : STD_LOGIC;
	signal p158_in : STD_LOGIC_VECTOR(0 to 91 - 1);
	signal p158_out : STD_LOGIC;
	signal p159_in : STD_LOGIC_VECTOR(0 to 105 - 1);
	signal p159_out : STD_LOGIC;
	signal p160_in : STD_LOGIC_VECTOR(0 to 178 - 1);
	signal p160_out : STD_LOGIC;
	signal p161_in : STD_LOGIC_VECTOR(0 to 85 - 1);
	signal p161_out : STD_LOGIC;
	signal p162_in : STD_LOGIC_VECTOR(0 to 83 - 1);
	signal p162_out : STD_LOGIC;
	signal p163_in : STD_LOGIC_VECTOR(0 to 107 - 1);
	signal p163_out : STD_LOGIC;
	signal p164_in : STD_LOGIC_VECTOR(0 to 84 - 1);
	signal p164_out : STD_LOGIC;
	signal p165_in : STD_LOGIC_VECTOR(0 to 166 - 1);
	signal p165_out : STD_LOGIC;
	signal p166_in : STD_LOGIC_VECTOR(0 to 129 - 1);
	signal p166_out : STD_LOGIC;
	signal p167_in : STD_LOGIC_VECTOR(0 to 90 - 1);
	signal p167_out : STD_LOGIC;
	signal p168_in : STD_LOGIC_VECTOR(0 to 176 - 1);
	signal p168_out : STD_LOGIC;
	signal p169_in : STD_LOGIC_VECTOR(0 to 131 - 1);
	signal p169_out : STD_LOGIC;
	signal p170_in : STD_LOGIC_VECTOR(0 to 110 - 1);
	signal p170_out : STD_LOGIC;
	signal p171_in : STD_LOGIC_VECTOR(0 to 95 - 1);
	signal p171_out : STD_LOGIC;
	signal p172_in : STD_LOGIC_VECTOR(0 to 248 - 1);
	signal p172_out : STD_LOGIC;
	signal p173_in : STD_LOGIC_VECTOR(0 to 107 - 1);
	signal p173_out : STD_LOGIC;
	signal p174_in : STD_LOGIC_VECTOR(0 to 165 - 1);
	signal p174_out : STD_LOGIC;
	signal p175_in : STD_LOGIC_VECTOR(0 to 138 - 1);
	signal p175_out : STD_LOGIC;
	signal p176_in : STD_LOGIC_VECTOR(0 to 49 - 1);
	signal p176_out : STD_LOGIC;
	signal p177_in : STD_LOGIC_VECTOR(0 to 151 - 1);
	signal p177_out : STD_LOGIC;
	signal p178_in : STD_LOGIC_VECTOR(0 to 108 - 1);
	signal p178_out : STD_LOGIC;
	signal p179_in : STD_LOGIC_VECTOR(0 to 101 - 1);
	signal p179_out : STD_LOGIC;
	signal p180_in : STD_LOGIC_VECTOR(0 to 114 - 1);
	signal p180_out : STD_LOGIC;
	signal p181_in : STD_LOGIC_VECTOR(0 to 82 - 1);
	signal p181_out : STD_LOGIC;
	signal p182_in : STD_LOGIC_VECTOR(0 to 104 - 1);
	signal p182_out : STD_LOGIC;
	signal p183_in : STD_LOGIC_VECTOR(0 to 74 - 1);
	signal p183_out : STD_LOGIC;
	signal p184_in : STD_LOGIC_VECTOR(0 to 97 - 1);
	signal p184_out : STD_LOGIC;
	signal p185_in : STD_LOGIC_VECTOR(0 to 118 - 1);
	signal p185_out : STD_LOGIC;
	signal p186_in : STD_LOGIC_VECTOR(0 to 152 - 1);
	signal p186_out : STD_LOGIC;
	signal p187_in : STD_LOGIC_VECTOR(0 to 91 - 1);
	signal p187_out : STD_LOGIC;
	signal p188_in : STD_LOGIC_VECTOR(0 to 120 - 1);
	signal p188_out : STD_LOGIC;
	signal p189_in : STD_LOGIC_VECTOR(0 to 100 - 1);
	signal p189_out : STD_LOGIC;
	signal p190_in : STD_LOGIC_VECTOR(0 to 68 - 1);
	signal p190_out : STD_LOGIC;
	signal p191_in : STD_LOGIC_VECTOR(0 to 90 - 1);
	signal p191_out : STD_LOGIC;
	signal p192_in : STD_LOGIC_VECTOR(0 to 64 - 1);
	signal p192_out : STD_LOGIC;
	signal p193_in : STD_LOGIC_VECTOR(0 to 118 - 1);
	signal p193_out : STD_LOGIC;
	signal p194_in : STD_LOGIC_VECTOR(0 to 66 - 1);
	signal p194_out : STD_LOGIC;
	signal p195_in : STD_LOGIC_VECTOR(0 to 74 - 1);
	signal p195_out : STD_LOGIC;
	signal p196_in : STD_LOGIC_VECTOR(0 to 97 - 1);
	signal p196_out : STD_LOGIC;
	signal p197_in : STD_LOGIC_VECTOR(0 to 116 - 1);
	signal p197_out : STD_LOGIC;
	signal p198_in : STD_LOGIC_VECTOR(0 to 194 - 1);
	signal p198_out : STD_LOGIC;
	signal p199_in : STD_LOGIC_VECTOR(0 to 115 - 1);
	signal p199_out : STD_LOGIC;
	signal p200_in : STD_LOGIC_VECTOR(0 to 253 - 1);
	signal p200_out : STD_LOGIC;
	signal p201_in : STD_LOGIC_VECTOR(0 to 89 - 1);
	signal p201_out : STD_LOGIC;
	signal p202_in : STD_LOGIC_VECTOR(0 to 132 - 1);
	signal p202_out : STD_LOGIC;
	signal p203_in : STD_LOGIC_VECTOR(0 to 112 - 1);
	signal p203_out : STD_LOGIC;
	signal p204_in : STD_LOGIC_VECTOR(0 to 138 - 1);
	signal p204_out : STD_LOGIC;
	signal p205_in : STD_LOGIC_VECTOR(0 to 74 - 1);
	signal p205_out : STD_LOGIC;
	signal p206_in : STD_LOGIC_VECTOR(0 to 99 - 1);
	signal p206_out : STD_LOGIC;
	signal p207_in : STD_LOGIC_VECTOR(0 to 78 - 1);
	signal p207_out : STD_LOGIC;
	signal p208_in : STD_LOGIC_VECTOR(0 to 114 - 1);
	signal p208_out : STD_LOGIC;
	signal p209_in : STD_LOGIC_VECTOR(0 to 111 - 1);
	signal p209_out : STD_LOGIC;
	signal p210_in : STD_LOGIC_VECTOR(0 to 104 - 1);
	signal p210_out : STD_LOGIC;
	signal p211_in : STD_LOGIC_VECTOR(0 to 60 - 1);
	signal p211_out : STD_LOGIC;
	signal p212_in : STD_LOGIC_VECTOR(0 to 78 - 1);
	signal p212_out : STD_LOGIC;
	signal p213_in : STD_LOGIC_VECTOR(0 to 69 - 1);
	signal p213_out : STD_LOGIC;
	signal p214_in : STD_LOGIC_VECTOR(0 to 92 - 1);
	signal p214_out : STD_LOGIC;
	signal p215_in : STD_LOGIC_VECTOR(0 to 92 - 1);
	signal p215_out : STD_LOGIC;
	signal p216_in : STD_LOGIC_VECTOR(0 to 122 - 1);
	signal p216_out : STD_LOGIC;
	signal p217_in : STD_LOGIC_VECTOR(0 to 72 - 1);
	signal p217_out : STD_LOGIC;
	signal p218_in : STD_LOGIC_VECTOR(0 to 133 - 1);
	signal p218_out : STD_LOGIC;
	signal p219_in : STD_LOGIC_VECTOR(0 to 89 - 1);
	signal p219_out : STD_LOGIC;
	signal p220_in : STD_LOGIC_VECTOR(0 to 73 - 1);
	signal p220_out : STD_LOGIC;
	signal p221_in : STD_LOGIC_VECTOR(0 to 115 - 1);
	signal p221_out : STD_LOGIC;
	signal p222_in : STD_LOGIC_VECTOR(0 to 114 - 1);
	signal p222_out : STD_LOGIC;
	signal p223_in : STD_LOGIC_VECTOR(0 to 73 - 1);
	signal p223_out : STD_LOGIC;
	signal p224_in : STD_LOGIC_VECTOR(0 to 102 - 1);
	signal p224_out : STD_LOGIC;
	signal p225_in : STD_LOGIC_VECTOR(0 to 64 - 1);
	signal p225_out : STD_LOGIC;
	signal p226_in : STD_LOGIC_VECTOR(0 to 145 - 1);
	signal p226_out : STD_LOGIC;
	signal p227_in : STD_LOGIC_VECTOR(0 to 117 - 1);
	signal p227_out : STD_LOGIC;
	signal p228_in : STD_LOGIC_VECTOR(0 to 65 - 1);
	signal p228_out : STD_LOGIC;
	signal p229_in : STD_LOGIC_VECTOR(0 to 119 - 1);
	signal p229_out : STD_LOGIC;
	signal p230_in : STD_LOGIC_VECTOR(0 to 57 - 1);
	signal p230_out : STD_LOGIC;
	signal p231_in : STD_LOGIC_VECTOR(0 to 187 - 1);
	signal p231_out : STD_LOGIC;
	signal p232_in : STD_LOGIC_VECTOR(0 to 48 - 1);
	signal p232_out : STD_LOGIC;
	signal p233_in : STD_LOGIC_VECTOR(0 to 86 - 1);
	signal p233_out : STD_LOGIC;
	signal p234_in : STD_LOGIC_VECTOR(0 to 104 - 1);
	signal p234_out : STD_LOGIC;
	signal p235_in : STD_LOGIC_VECTOR(0 to 127 - 1);
	signal p235_out : STD_LOGIC;
	signal p236_in : STD_LOGIC_VECTOR(0 to 78 - 1);
	signal p236_out : STD_LOGIC;
	signal p237_in : STD_LOGIC_VECTOR(0 to 101 - 1);
	signal p237_out : STD_LOGIC;
	signal p238_in : STD_LOGIC_VECTOR(0 to 76 - 1);
	signal p238_out : STD_LOGIC;
	signal p239_in : STD_LOGIC_VECTOR(0 to 136 - 1);
	signal p239_out : STD_LOGIC;
	signal p240_in : STD_LOGIC_VECTOR(0 to 103 - 1);
	signal p240_out : STD_LOGIC;
	signal p241_in : STD_LOGIC_VECTOR(0 to 132 - 1);
	signal p241_out : STD_LOGIC;
	signal p242_in : STD_LOGIC_VECTOR(0 to 78 - 1);
	signal p242_out : STD_LOGIC;
	signal p243_in : STD_LOGIC_VECTOR(0 to 85 - 1);
	signal p243_out : STD_LOGIC;
	signal p244_in : STD_LOGIC_VECTOR(0 to 218 - 1);
	signal p244_out : STD_LOGIC;
	signal p245_in : STD_LOGIC_VECTOR(0 to 119 - 1);
	signal p245_out : STD_LOGIC;
	signal p246_in : STD_LOGIC_VECTOR(0 to 98 - 1);
	signal p246_out : STD_LOGIC;
	signal p247_in : STD_LOGIC_VECTOR(0 to 61 - 1);
	signal p247_out : STD_LOGIC;
	signal p248_in : STD_LOGIC_VECTOR(0 to 119 - 1);
	signal p248_out : STD_LOGIC;
	signal p249_in : STD_LOGIC_VECTOR(0 to 82 - 1);
	signal p249_out : STD_LOGIC;
	signal p250_in : STD_LOGIC_VECTOR(0 to 119 - 1);
	signal p250_out : STD_LOGIC;
	signal p251_in : STD_LOGIC_VECTOR(0 to 107 - 1);
	signal p251_out : STD_LOGIC;
	signal p252_in : STD_LOGIC_VECTOR(0 to 106 - 1);
	signal p252_out : STD_LOGIC;
	signal p253_in : STD_LOGIC_VECTOR(0 to 129 - 1);
	signal p253_out : STD_LOGIC;
	signal p254_in : STD_LOGIC_VECTOR(0 to 127 - 1);
	signal p254_out : STD_LOGIC;
	signal p255_in : STD_LOGIC_VECTOR(0 to 90 - 1);
	signal p255_out : STD_LOGIC;
	
    
    -- Dummies
    signal dummy0 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy1 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy2 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy3 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy4 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy5 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy6 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy7 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy8 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy9 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy10 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy11 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy12 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy13 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy14 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy15 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy16 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy17 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy18 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy19 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy20 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy21 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy22 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy23 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy24 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy25 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy26 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy27 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy28 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy29 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy30 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy31 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy32 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy33 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy34 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy35 : STD_LOGIC_VECTOR(0 to 18 - 2);
	signal dummy36 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy37 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy38 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy39 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy40 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy41 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy42 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy43 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy44 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy45 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy46 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy47 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy48 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy49 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy50 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy51 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy52 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy53 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy54 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy55 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy56 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy57 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy58 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy59 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy60 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy61 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy62 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy63 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy64 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy65 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy66 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy67 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy68 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy69 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy70 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy71 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy72 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy73 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy74 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy75 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy76 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy77 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy78 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy79 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy80 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy81 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy82 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy83 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy84 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy85 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy86 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy87 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy88 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy89 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy90 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy91 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy92 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy93 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy94 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy95 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy96 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy97 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy98 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy99 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy100 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy101 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy102 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy103 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy104 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy105 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy106 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy107 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy108 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy109 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy110 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy111 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy112 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy113 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy114 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy115 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy116 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy117 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy118 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy119 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy120 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy121 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy122 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy123 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy124 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy125 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy126 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy127 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy128 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy129 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy130 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy131 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy132 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy133 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy134 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy135 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy136 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy137 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy138 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy139 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy140 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy141 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy142 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy143 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy144 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy145 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy146 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy147 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy148 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy149 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy150 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy151 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy152 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy153 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy154 : STD_LOGIC_VECTOR(0 to 18 - 2);
	signal dummy155 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy156 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy157 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy158 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy159 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy160 : STD_LOGIC_VECTOR(0 to 18 - 2);
	signal dummy161 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy162 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy163 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy164 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy165 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy166 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy167 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy168 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy169 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy170 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy171 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy172 : STD_LOGIC_VECTOR(0 to 18 - 2);
	signal dummy173 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy174 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy175 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy176 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy177 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy178 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy179 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy180 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy181 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy182 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy183 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy184 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy185 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy186 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy187 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy188 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy189 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy190 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy191 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy192 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy193 : STD_LOGIC_VECTOR(0 to 18 - 2);
	signal dummy194 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy195 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy196 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy197 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy198 : STD_LOGIC_VECTOR(0 to 18 - 2);
	signal dummy199 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy200 : STD_LOGIC_VECTOR(0 to 18 - 2);
	signal dummy201 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy202 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy203 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy204 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy205 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy206 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy207 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy208 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy209 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy210 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy211 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy212 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy213 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy214 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy215 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy216 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy217 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy218 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy219 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy220 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy221 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy222 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy223 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy224 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy225 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy226 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy227 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy228 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy229 : STD_LOGIC_VECTOR(0 to 18 - 2);
	signal dummy230 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy231 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy232 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy233 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy234 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy235 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy236 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy237 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy238 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy239 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy240 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy241 : STD_LOGIC_VECTOR(0 to 18 - 2);
	signal dummy242 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy243 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy244 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy245 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy246 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy247 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy248 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy249 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy250 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy251 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy252 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy253 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy254 : STD_LOGIC_VECTOR(0 to 17 - 2);
	signal dummy255 : STD_LOGIC_VECTOR(0 to 16 - 2);
	 

begin

    
    p0_in <= x(101) & x(102) & x(103) & x(200) & x(220) & x(221) & x(227) & x(247) & x(248) & x(249) & x(250) & x(275) & x(276) & x(277) & x(278) & x(297) & x(306) & x(324) & x(325) & x(348) & x(349) & x(350) & x(377) & x(378) & x(405) & x(406) & x(433) & x(436) & x(464) & x(542) & x(570) & x(708) & x(735) & x(737) & x(738) & x(739);
    y(0) <= not(p0_out);
    p0 : perceptron
        Generic map (
            WEIGHTS => "111100100000000101100000000110011111",
            SHIFT => 4,
            B => -56,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p0_in,
            y(0) => p0_out,
            y(1 to 15 - 1) => dummy0
        );


    p1_in <= x(70) & x(72) & x(73) & x(75) & x(78) & x(104) & x(105) & x(154) & x(155) & x(157) & x(198) & x(199) & x(201) & x(203) & x(226) & x(227) & x(241) & x(249) & x(250) & x(254) & x(255) & x(267) & x(268) & x(269) & x(282) & x(283) & x(284) & x(294) & x(295) & x(309) & x(310) & x(311) & x(312) & x(317) & x(318) & x(319) & x(322) & x(323) & x(338) & x(339) & x(345) & x(353) & x(355) & x(356) & x(361) & x(362) & x(366) & x(367) & x(372) & x(373) & x(376) & x(377) & x(378) & x(381) & x(383) & x(404) & x(405) & x(406) & x(409) & x(432) & x(433) & x(436) & x(457) & x(458) & x(459) & x(460) & x(461) & x(464) & x(487) & x(488) & x(508) & x(514) & x(515) & x(535) & x(536) & x(564) & x(571) & x(592) & x(593) & x(599) & x(620) & x(624) & x(625) & x(648) & x(649) & x(653) & x(654) & x(666) & x(677) & x(678) & x(693) & x(694) & x(695) & x(696) & x(704) & x(706) & x(707) & x(708) & x(719) & x(720) & x(721) & x(722) & x(723) & x(735) & x(736) & x(743) & x(748) & x(749) & x(764) & x(765) & x(766) & x(769) & x(770) & x(771) & x(772) & x(773) & x(774);
    y(1) <= not(p1_out);
    p1 : perceptron
        Generic map (
            WEIGHTS => "000000011111111111111111111111111000111100001111000000000000000000000010011111111111111011000011110000011100111111111",
            SHIFT => 3,
            B => 293,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p1_in,
            y(0) => p1_out,
            y(1 to 16 - 1) => dummy1
        );


    p2_in <= x(34) & x(37) & x(40) & x(41) & x(62) & x(63) & x(64) & x(65) & x(66) & x(118) & x(122) & x(154) & x(155) & x(198) & x(199) & x(202) & x(226) & x(227) & x(228) & x(237) & x(248) & x(249) & x(254) & x(255) & x(256) & x(266) & x(267) & x(268) & x(276) & x(277) & x(282) & x(283) & x(284) & x(294) & x(295) & x(296) & x(297) & x(309) & x(310) & x(311) & x(312) & x(316) & x(318) & x(320) & x(337) & x(338) & x(339) & x(342) & x(345) & x(346) & x(347) & x(348) & x(349) & x(353) & x(362) & x(366) & x(367) & x(370) & x(371) & x(372) & x(378) & x(379) & x(381) & x(387) & x(390) & x(396) & x(398) & x(409) & x(418) & x(424) & x(430) & x(431) & x(433) & x(436) & x(446) & x(458) & x(459) & x(468) & x(473) & x(474) & x(481) & x(487) & x(495) & x(497) & x(500) & x(501) & x(502) & x(509) & x(528) & x(529) & x(530) & x(555) & x(556) & x(557) & x(558) & x(564) & x(569) & x(583) & x(584) & x(585) & x(599) & x(611) & x(612) & x(638) & x(640) & x(690) & x(691) & x(692) & x(693) & x(694) & x(695) & x(696) & x(706) & x(707) & x(708) & x(719) & x(720) & x(721) & x(722) & x(723) & x(735) & x(736) & x(737) & x(741) & x(742) & x(743) & x(744) & x(748) & x(749) & x(764) & x(765) & x(766) & x(769) & x(770) & x(771) & x(772) & x(773) & x(774);
    y(2) <= not(p2_out);
    p2 : perceptron
        Generic map (
            WEIGHTS => "000000000111111111110011111100111111111110001110000000111000000010001000001001111011111111111111111111111000000011100000111111100111111111",
            SHIFT => 4,
            B => 482,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p2_in,
            y(0) => p2_out,
            y(1 to 17 - 1) => dummy2
        );


    p3_in <= x(65) & x(66) & x(102) & x(103) & x(108) & x(118) & x(135) & x(163) & x(164) & x(165) & x(166) & x(191) & x(192) & x(193) & x(194) & x(215) & x(219) & x(220) & x(221) & x(222) & x(239) & x(247) & x(248) & x(249) & x(250) & x(273) & x(276) & x(277) & x(278) & x(295) & x(297) & x(303) & x(305) & x(309) & x(328) & x(329) & x(330) & x(331) & x(332) & x(338) & x(342) & x(347) & x(348) & x(350) & x(368) & x(370) & x(375) & x(376) & x(377) & x(390) & x(418) & x(446) & x(473) & x(474) & x(481) & x(501) & x(502) & x(529) & x(544) & x(545) & x(557) & x(558) & x(584) & x(640) & x(652) & x(655) & x(656) & x(657) & x(658) & x(693) & x(694);
    y(3) <= not(p3_out);
    p3 : perceptron
        Generic map (
            WEIGHTS => "11000011111111111111011111111000100000001111111110000000000000001111111",
            SHIFT => 4,
            B => 104,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p3_in,
            y(0) => p3_out,
            y(1 to 16 - 1) => dummy3
        );


    p4_in <= x(37) & x(65) & x(93) & x(94) & x(95) & x(96) & x(97) & x(98) & x(99) & x(104) & x(105) & x(123) & x(124) & x(125) & x(126) & x(127) & x(138) & x(153) & x(162) & x(163) & x(166) & x(182) & x(183) & x(184) & x(190) & x(191) & x(210) & x(211) & x(212) & x(233) & x(238) & x(239) & x(248) & x(249) & x(250) & x(276) & x(277) & x(304) & x(306) & x(311) & x(334) & x(346) & x(387) & x(390) & x(418) & x(422) & x(438) & x(439) & x(444) & x(446) & x(463) & x(471) & x(474) & x(487) & x(498) & x(499) & x(500) & x(501) & x(502) & x(514) & x(528) & x(529) & x(541) & x(542) & x(556) & x(557) & x(583) & x(584) & x(622) & x(694) & x(695) & x(712) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(732) & x(742) & x(745) & x(746) & x(747) & x(748) & x(749) & x(769) & x(771);
    y(4) <= not(p4_out);
    p4 : perceptron
        Generic map (
            WEIGHTS => "01111111100111111100111100111011111111101001100011011111111111111111111111111111111111100",
            SHIFT => 4,
            B => 848,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p4_in,
            y(0) => p4_out,
            y(1 to 16 - 1) => dummy4
        );


    p5_in <= x(67) & x(68) & x(69) & x(91) & x(108) & x(151) & x(152) & x(182) & x(184) & x(191) & x(192) & x(209) & x(210) & x(211) & x(212) & x(213) & x(238) & x(239) & x(305) & x(307) & x(333) & x(334) & x(361) & x(362) & x(433) & x(462) & x(463) & x(490) & x(529) & x(594) & x(622) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(732) & x(739) & x(742) & x(744) & x(745) & x(746) & x(747) & x(748) & x(749);
    y(5) <= not(p5_out);
    p5 : perceptron
        Generic map (
            WEIGHTS => "11111111100111111100000000001111111111111111111",
            SHIFT => 4,
            B => 346,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p5_in,
            y(0) => p5_out,
            y(1 to 15 - 1) => dummy5
        );


    p6_in <= x(68) & x(70) & x(74) & x(75) & x(77) & x(78) & x(79) & x(101) & x(102) & x(103) & x(104) & x(105) & x(106) & x(107) & x(108) & x(166) & x(182) & x(187) & x(188) & x(192) & x(193) & x(194) & x(198) & x(221) & x(222) & x(227) & x(228) & x(248) & x(249) & x(250) & x(254) & x(264) & x(265) & x(268) & x(276) & x(277) & x(278) & x(283) & x(296) & x(297) & x(299) & x(300) & x(302) & x(305) & x(306) & x(309) & x(310) & x(311) & x(326) & x(327) & x(328) & x(329) & x(330) & x(331) & x(332) & x(333) & x(334) & x(337) & x(338) & x(339) & x(349) & x(350) & x(357) & x(358) & x(359) & x(360) & x(362) & x(366) & x(377) & x(378) & x(387) & x(394) & x(406) & x(418) & x(461) & x(485) & x(513) & x(514) & x(515) & x(550) & x(595) & x(596) & x(620) & x(624) & x(646) & x(707) & x(711) & x(712) & x(713) & x(714) & x(719) & x(720) & x(721) & x(723) & x(735) & x(738) & x(742) & x(743) & x(769) & x(770) & x(771) & x(772) & x(773) & x(774);
    y(6) <= not(p6_out);
    p6 : perceptron
        Generic map (
            WEIGHTS => "00000000000000011111110110011100001110000001100000000001100011000010110011100001111110000011110000000000",
            SHIFT => 4,
            B => -402,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p6_in,
            y(0) => p6_out,
            y(1 to 16 - 1) => dummy6
        );


    p7_in <= x(34) & x(35) & x(36) & x(37) & x(38) & x(39) & x(40) & x(41) & x(42) & x(44) & x(45) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(79) & x(80) & x(90) & x(91) & x(92) & x(93) & x(94) & x(95) & x(96) & x(97) & x(98) & x(99) & x(100) & x(101) & x(102) & x(103) & x(104) & x(105) & x(106) & x(107) & x(108) & x(135) & x(162) & x(163) & x(164) & x(186) & x(192) & x(277) & x(303) & x(304) & x(323) & x(330) & x(331) & x(332) & x(338) & x(353) & x(358) & x(359) & x(368) & x(382) & x(387) & x(388) & x(397) & x(401) & x(436) & x(464) & x(514) & x(515) & x(516) & x(541) & x(542) & x(543) & x(544) & x(571) & x(693) & x(694) & x(719);
    y(7) <= not(p7_out);
    p7 : perceptron
        Generic map (
            WEIGHTS => "0000000000000000000000000000000000000000000000000111111100100000001000110000000000111",
            SHIFT => 4,
            B => -904,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p7_in,
            y(0) => p7_out,
            y(1 to 16 - 1) => dummy7
        );


    p8_in <= x(152) & x(153) & x(154) & x(155) & x(181) & x(192) & x(220) & x(221) & x(222) & x(248) & x(249) & x(250) & x(276) & x(277) & x(278) & x(330) & x(358) & x(373) & x(374) & x(378) & x(400) & x(402) & x(405) & x(406) & x(432) & x(433) & x(434) & x(440) & x(441) & x(473) & x(501) & x(514) & x(515) & x(516) & x(675) & x(677) & x(678) & x(705) & x(706) & x(707) & x(708) & x(709);
    y(8) <= not(p8_out);
    p8 : perceptron
        Generic map (
            WEIGHTS => "000001111111111001101100000110000011111111",
            SHIFT => 4,
            B => 247,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p8_in,
            y(0) => p8_out,
            y(1 to 15 - 1) => dummy8
        );


    p9_in <= x(74) & x(75) & x(76) & x(103) & x(104) & x(106) & x(107) & x(108) & x(198) & x(210) & x(221) & x(222) & x(233) & x(238) & x(239) & x(249) & x(267) & x(277) & x(289) & x(292) & x(295) & x(309) & x(320) & x(330) & x(331) & x(343) & x(344) & x(347) & x(348) & x(350) & x(353) & x(357) & x(359) & x(361) & x(403) & x(408) & x(431) & x(436) & x(473) & x(474) & x(479) & x(485) & x(501) & x(502) & x(507) & x(513) & x(514) & x(515) & x(528) & x(529) & x(530) & x(535) & x(556) & x(557) & x(558) & x(563) & x(583) & x(584) & x(585) & x(591) & x(592) & x(611) & x(612) & x(619) & x(620) & x(636) & x(637) & x(638) & x(640) & x(666) & x(691) & x(692) & x(716) & x(743) & x(773);
    y(9) <= not(p9_out);
    p9 : perceptron
        Generic map (
            WEIGHTS => "111111111000100000110111111110111111110001000111000000000000000000000011111",
            SHIFT => 4,
            B => -126,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p9_in,
            y(0) => p9_out,
            y(1 to 16 - 1) => dummy9
        );


    p10_in <= x(34) & x(35) & x(37) & x(38) & x(39) & x(40) & x(41) & x(62) & x(63) & x(64) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(78) & x(79) & x(95) & x(96) & x(97) & x(100) & x(101) & x(102) & x(103) & x(104) & x(105) & x(136) & x(165) & x(166) & x(192) & x(193) & x(198) & x(220) & x(221) & x(247) & x(248) & x(249) & x(250) & x(262) & x(263) & x(274) & x(275) & x(276) & x(277) & x(278) & x(289) & x(290) & x(291) & x(304) & x(305) & x(306) & x(307) & x(319) & x(320) & x(333) & x(334) & x(341) & x(347) & x(348) & x(349) & x(358) & x(359) & x(360) & x(362) & x(368) & x(376) & x(386) & x(387) & x(388) & x(418) & x(446) & x(543) & x(591) & x(619) & x(692) & x(711) & x(712) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(744) & x(745) & x(746) & x(747) & x(748) & x(773);
    y(10) <= not(p10_out);
    p10 : perceptron
        Generic map (
            WEIGHTS => "111111111111111111111111111111100000000000000000000000000000000001110001110011100000000000000000",
            SHIFT => 4,
            B => -197,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p10_in,
            y(0) => p10_out,
            y(1 to 16 - 1) => dummy10
        );


    p11_in <= x(64) & x(108) & x(118) & x(124) & x(125) & x(126) & x(135) & x(162) & x(163) & x(164) & x(165) & x(171) & x(172) & x(181) & x(182) & x(188) & x(189) & x(190) & x(191) & x(192) & x(193) & x(194) & x(200) & x(210) & x(211) & x(217) & x(218) & x(219) & x(220) & x(221) & x(222) & x(226) & x(238) & x(239) & x(247) & x(248) & x(249) & x(250) & x(260) & x(263) & x(276) & x(277) & x(288) & x(289) & x(291) & x(296) & x(303) & x(304) & x(316) & x(320) & x(327) & x(328) & x(329) & x(330) & x(331) & x(332) & x(343) & x(345) & x(346) & x(347) & x(348) & x(360) & x(390) & x(397) & x(398) & x(418) & x(425) & x(446) & x(450) & x(474) & x(475) & x(479) & x(502) & x(507) & x(534) & x(535) & x(557) & x(562) & x(563) & x(591) & x(618) & x(619) & x(620) & x(646) & x(647) & x(648) & x(668) & x(694) & x(695) & x(704) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(745) & x(746) & x(747) & x(748) & x(749);
    y(11) <= not(p11_out);
    p11 : perceptron
        Generic map (
            WEIGHTS => "1000001111100001111111000111111100111111111110001100000011111001101000000000000000000000010000000000000",
            SHIFT => 4,
            B => -352,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p11_in,
            y(0) => p11_out,
            y(1 to 16 - 1) => dummy11
        );


    p12_in <= x(40) & x(46) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(103) & x(131) & x(132) & x(156) & x(157) & x(175) & x(202) & x(204) & x(221) & x(222) & x(230) & x(231) & x(248) & x(249) & x(250) & x(276) & x(277) & x(292) & x(297) & x(299) & x(302) & x(303) & x(311) & x(326) & x(329) & x(330) & x(337) & x(339) & x(341) & x(342) & x(369) & x(370) & x(371) & x(374) & x(386) & x(413) & x(414) & x(433) & x(442) & x(444) & x(469) & x(473) & x(474) & x(491) & x(501) & x(502) & x(514) & x(528) & x(529) & x(530) & x(556) & x(557) & x(558) & x(572) & x(582) & x(583) & x(584) & x(609) & x(610) & x(611) & x(612) & x(634) & x(635) & x(636) & x(637) & x(638) & x(675) & x(677) & x(678) & x(694) & x(695) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(747) & x(748) & x(749) & x(773) & x(774);
    y(12) <= not(p12_out);
    p12 : perceptron
        Generic map (
            WEIGHTS => "0000000000000001111100110000001111111111000000000100011111111111101111111111110000000000000011",
            SHIFT => 4,
            B => -205,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p12_in,
            y(0) => p12_out,
            y(1 to 16 - 1) => dummy12
        );


    p13_in <= x(78) & x(79) & x(104) & x(105) & x(106) & x(164) & x(165) & x(166) & x(192) & x(193) & x(194) & x(220) & x(221) & x(222) & x(247) & x(248) & x(249) & x(250) & x(275) & x(276) & x(277) & x(278) & x(304) & x(305) & x(306) & x(321) & x(322) & x(333) & x(334) & x(348) & x(349) & x(350) & x(358) & x(359) & x(360) & x(361) & x(362) & x(377) & x(378) & x(385) & x(386) & x(387) & x(388) & x(390) & x(425) & x(426) & x(453) & x(454) & x(501) & x(529) & x(557) & x(558) & x(584) & x(612) & x(656) & x(657) & x(720) & x(721) & x(764);
    y(13) <= not(p13_out);
    p13 : perceptron
        Generic map (
            WEIGHTS => "11111000000000000000000000000000111000011110111111111100000",
            SHIFT => 4,
            B => -210,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p13_in,
            y(0) => p13_out,
            y(1 to 16 - 1) => dummy13
        );


    p14_in <= x(35) & x(39) & x(40) & x(41) & x(43) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(101) & x(102) & x(103) & x(104) & x(105) & x(106) & x(158) & x(187) & x(188) & x(217) & x(233) & x(234) & x(242) & x(246) & x(247) & x(249) & x(261) & x(266) & x(267) & x(276) & x(277) & x(297) & x(298) & x(299) & x(301) & x(302) & x(303) & x(329) & x(330) & x(331) & x(332) & x(333) & x(338) & x(352) & x(353) & x(361) & x(372) & x(375) & x(376) & x(380) & x(381) & x(384) & x(387) & x(388) & x(398) & x(399) & x(400) & x(402) & x(403) & x(404) & x(408) & x(412) & x(414) & x(415) & x(416) & x(418) & x(427) & x(430) & x(431) & x(433) & x(436) & x(437) & x(444) & x(446) & x(473) & x(474) & x(475) & x(501) & x(502) & x(515) & x(529) & x(530) & x(549) & x(557) & x(558) & x(576) & x(582) & x(583) & x(584) & x(598) & x(612) & x(640) & x(657) & x(659) & x(660) & x(703) & x(704) & x(737) & x(739) & x(742) & x(743) & x(745) & x(746) & x(770) & x(772);
    y(14) <= not(p14_out);
    p14 : perceptron
        Generic map (
            WEIGHTS => "111111111111111111111111111100000000010001100000000000011011111111111111111110111011100000000010010000000001100000000",
            SHIFT => 4,
            B => 25,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p14_in,
            y(0) => p14_out,
            y(1 to 17 - 1) => dummy14
        );


    p15_in <= x(63) & x(79) & x(96) & x(108) & x(126) & x(127) & x(134) & x(135) & x(136) & x(154) & x(155) & x(156) & x(161) & x(162) & x(163) & x(164) & x(165) & x(166) & x(184) & x(191) & x(192) & x(193) & x(194) & x(219) & x(220) & x(221) & x(222) & x(247) & x(248) & x(249) & x(250) & x(251) & x(276) & x(277) & x(278) & x(298) & x(300) & x(302) & x(303) & x(305) & x(306) & x(307) & x(322) & x(323) & x(328) & x(329) & x(330) & x(331) & x(332) & x(333) & x(334) & x(338) & x(342) & x(349) & x(350) & x(357) & x(358) & x(359) & x(360) & x(361) & x(362) & x(370) & x(371) & x(373) & x(378) & x(399) & x(450) & x(454) & x(473) & x(474) & x(478) & x(481) & x(483) & x(485) & x(501) & x(502) & x(506) & x(507) & x(512) & x(513) & x(514) & x(515) & x(529) & x(530) & x(535) & x(542) & x(543) & x(556) & x(557) & x(558) & x(584) & x(612) & x(638) & x(640) & x(648) & x(675) & x(676) & x(677) & x(678) & x(679) & x(732) & x(745) & x(746) & x(747);
    y(15) <= not(p15_out);
    p15 : perceptron
        Generic map (
            WEIGHTS => "00000011100011111101111111111111111000011111000001101110000111111110001000001100000010000000001111110000",
            SHIFT => 4,
            B => 103,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p15_in,
            y(0) => p15_out,
            y(1 to 16 - 1) => dummy15
        );


    p16_in <= x(35) & x(44) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(70) & x(75) & x(76) & x(91) & x(92) & x(93) & x(94) & x(95) & x(96) & x(101) & x(102) & x(103) & x(104) & x(148) & x(156) & x(163) & x(182) & x(198) & x(199) & x(227) & x(242) & x(248) & x(249) & x(250) & x(269) & x(276) & x(277) & x(295) & x(306) & x(322) & x(325) & x(370) & x(386) & x(410) & x(414) & x(431) & x(437) & x(458) & x(459) & x(473) & x(474) & x(486) & x(487) & x(500) & x(501) & x(502) & x(512) & x(514) & x(528) & x(529) & x(540) & x(541) & x(542) & x(543) & x(555) & x(556) & x(557) & x(570) & x(575) & x(583) & x(584) & x(610) & x(611) & x(612) & x(638) & x(640) & x(693) & x(694) & x(706) & x(707) & x(708) & x(735) & x(736) & x(737) & x(743) & x(746);
    y(16) <= not(p16_out);
    p16 : perceptron
        Generic map (
            WEIGHTS => "111111111111111111111010100001110110100010110111111111111111111111111111110000000000",
            SHIFT => 4,
            B => 514,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p16_in,
            y(0) => p16_out,
            y(1 to 16 - 1) => dummy16
        );


    p17_in <= x(34) & x(35) & x(36) & x(37) & x(38) & x(39) & x(40) & x(63) & x(66) & x(68) & x(117) & x(171) & x(172) & x(173) & x(200) & x(219) & x(247) & x(248) & x(275) & x(290) & x(291) & x(292) & x(295) & x(303) & x(305) & x(317) & x(319) & x(323) & x(330) & x(333) & x(418) & x(450) & x(473) & x(474) & x(479) & x(501) & x(502) & x(507) & x(515) & x(524) & x(528) & x(529) & x(530) & x(534) & x(535) & x(552) & x(556) & x(557) & x(558) & x(563) & x(570) & x(571) & x(584) & x(585) & x(591) & x(592) & x(612) & x(618) & x(619) & x(620) & x(647) & x(648) & x(649) & x(658) & x(675) & x(676) & x(677) & x(678);
    y(17) <= not(p17_out);
    p17 : perceptron
        Generic map (
            WEIGHTS => "11111111110000011111110101101000000000100000000000000000000000010000",
            SHIFT => 5,
            B => -613,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p17_in,
            y(0) => p17_out,
            y(1 to 17 - 1) => dummy17
        );


    p18_in <= x(37) & x(38) & x(39) & x(40) & x(41) & x(45) & x(46) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(79) & x(102) & x(103) & x(104) & x(105) & x(108) & x(152) & x(163) & x(183) & x(192) & x(198) & x(208) & x(210) & x(211) & x(226) & x(235) & x(236) & x(239) & x(263) & x(264) & x(275) & x(277) & x(301) & x(302) & x(303) & x(304) & x(305) & x(328) & x(329) & x(330) & x(331) & x(332) & x(353) & x(354) & x(361) & x(362) & x(366) & x(381) & x(389) & x(390) & x(394) & x(397) & x(398) & x(400) & x(402) & x(413) & x(414) & x(418) & x(425) & x(426) & x(427) & x(440) & x(446) & x(450) & x(474) & x(507) & x(514) & x(535) & x(563) & x(573) & x(591) & x(602) & x(648) & x(649) & x(675) & x(676) & x(677) & x(678) & x(690) & x(691) & x(692) & x(703) & x(709) & x(711) & x(712) & x(713) & x(714) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(736) & x(737) & x(740) & x(741) & x(742) & x(744) & x(745) & x(746) & x(747) & x(748) & x(750) & x(771) & x(772);
    y(18) <= not(p18_out);
    p18 : perceptron
        Generic map (
            WEIGHTS => "1111111111111111111111111111100101000000000001000010000000000000011111101111010101111111111100010000000000000000000000000",
            SHIFT => 4,
            B => 47,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p18_in,
            y(0) => p18_out,
            y(1 to 17 - 1) => dummy18
        );


    p19_in <= x(41) & x(69) & x(71) & x(72) & x(73) & x(74) & x(75) & x(93) & x(163) & x(192) & x(194) & x(221) & x(222) & x(248) & x(249) & x(250) & x(276) & x(277) & x(278) & x(302) & x(303) & x(304) & x(305) & x(306) & x(309) & x(320) & x(321) & x(322) & x(323) & x(329) & x(330) & x(331) & x(332) & x(348) & x(357) & x(358) & x(359) & x(360) & x(361) & x(368) & x(386) & x(387) & x(388) & x(414) & x(416) & x(443) & x(444) & x(446) & x(451) & x(468) & x(473) & x(474) & x(479) & x(489) & x(501) & x(502) & x(507) & x(518) & x(528) & x(529) & x(530) & x(534) & x(556) & x(557) & x(584) & x(611) & x(612) & x(628) & x(629) & x(636) & x(637) & x(638) & x(657) & x(660) & x(666) & x(682) & x(683) & x(693) & x(694) & x(710) & x(712) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(732) & x(747) & x(748) & x(749);
    y(19) <= not(p19_out);
    p19 : perceptron
        Generic map (
            WEIGHTS => "11111110000000000001110011100111111111101111111001000000000001000001100011011000000000000000",
            SHIFT => 4,
            B => -413,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p19_in,
            y(0) => p19_out,
            y(1 to 16 - 1) => dummy19
        );


    p20_in <= x(35) & x(37) & x(38) & x(40) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(79) & x(91) & x(96) & x(97) & x(98) & x(99) & x(100) & x(101) & x(102) & x(103) & x(104) & x(105) & x(106) & x(107) & x(108) & x(135) & x(136) & x(163) & x(164) & x(165) & x(166) & x(181) & x(182) & x(183) & x(184) & x(190) & x(191) & x(192) & x(193) & x(209) & x(210) & x(211) & x(212) & x(218) & x(219) & x(220) & x(221) & x(222) & x(237) & x(238) & x(239) & x(247) & x(248) & x(249) & x(266) & x(276) & x(277) & x(302) & x(305) & x(320) & x(328) & x(329) & x(330) & x(331) & x(332) & x(334) & x(347) & x(348) & x(357) & x(358) & x(359) & x(386) & x(387) & x(450) & x(487) & x(513) & x(514) & x(515) & x(516) & x(535) & x(542) & x(543) & x(647) & x(675) & x(676) & x(694) & x(695) & x(703) & x(712) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(732) & x(738) & x(739) & x(740) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(748) & x(749) & x(769);
    y(20) <= not(p20_out);
    p20 : perceptron
        Generic map (
            WEIGHTS => "1111111111111111111111111111111111100000011110000111100000111000100100111110001111101111101100011011111111111111111111110",
            SHIFT => 4,
            B => 565,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p20_in,
            y(0) => p20_out,
            y(1 to 17 - 1) => dummy20
        );


    p21_in <= x(166) & x(193) & x(198) & x(219) & x(220) & x(221) & x(247) & x(248) & x(249) & x(250) & x(255) & x(261) & x(262) & x(275) & x(276) & x(277) & x(278) & x(288) & x(289) & x(290) & x(303) & x(304) & x(305) & x(306) & x(307) & x(316) & x(319) & x(320) & x(333) & x(334) & x(347) & x(348) & x(349) & x(361) & x(362) & x(375) & x(376) & x(377) & x(390) & x(413) & x(414) & x(441) & x(442) & x(450) & x(470) & x(498) & x(510) & x(526) & x(537) & x(541) & x(557) & x(564) & x(565) & x(592) & x(620) & x(621) & x(655) & x(656) & x(657) & x(658) & x(685) & x(739) & x(746);
    y(21) <= not(p21_out);
    p21 : perceptron
        Generic map (
            WEIGHTS => "001000000000000000000000000000000000000111101111101111110000011",
            SHIFT => 4,
            B => -287,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p21_in,
            y(0) => p21_out,
            y(1 to 16 - 1) => dummy21
        );


    p22_in <= x(35) & x(62) & x(63) & x(64) & x(67) & x(68) & x(105) & x(108) & x(164) & x(165) & x(166) & x(191) & x(192) & x(193) & x(194) & x(198) & x(216) & x(217) & x(220) & x(221) & x(222) & x(226) & x(246) & x(248) & x(249) & x(250) & x(251) & x(266) & x(267) & x(276) & x(277) & x(278) & x(293) & x(294) & x(295) & x(298) & x(305) & x(306) & x(309) & x(310) & x(333) & x(334) & x(338) & x(339) & x(347) & x(348) & x(349) & x(350) & x(357) & x(358) & x(359) & x(366) & x(376) & x(377) & x(378) & x(386) & x(404) & x(432) & x(433) & x(450) & x(460) & x(461) & x(479) & x(488) & x(507) & x(535) & x(591) & x(647) & x(675) & x(736) & x(739) & x(741) & x(742) & x(743) & x(744) & x(746) & x(764) & x(770) & x(773) & x(774);
    y(22) <= not(p22_out);
    p22 : perceptron
        Generic map (
            WEIGHTS => "11111111000000010000010000011000111100110011000011110001000000000000011111111111",
            SHIFT => 4,
            B => -52,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p22_in,
            y(0) => p22_out,
            y(1 to 16 - 1) => dummy22
        );


    p23_in <= x(0) & x(8) & x(11) & x(22) & x(23) & x(52) & x(53) & x(54) & x(55) & x(56) & x(66) & x(71) & x(88) & x(98) & x(99) & x(108) & x(111) & x(113) & x(141) & x(153) & x(154) & x(155) & x(165) & x(167) & x(168) & x(169) & x(171) & x(181) & x(182) & x(196) & x(197) & x(199) & x(200) & x(220) & x(221) & x(222) & x(227) & x(248) & x(249) & x(250) & x(254) & x(255) & x(277) & x(283) & x(294) & x(295) & x(339) & x(364) & x(366) & x(370) & x(371) & x(372) & x(373) & x(392) & x(398) & x(399) & x(400) & x(401) & x(405) & x(406) & x(428) & x(432) & x(433) & x(440) & x(441) & x(442) & x(450) & x(453) & x(460) & x(461) & x(467) & x(468) & x(473) & x(483) & x(487) & x(488) & x(501) & x(503) & x(512) & x(513) & x(514) & x(515) & x(516) & x(518) & x(528) & x(529) & x(530) & x(557) & x(558) & x(560) & x(584) & x(612) & x(617) & x(636) & x(640) & x(667) & x(675) & x(676) & x(677) & x(678) & x(679) & x(701) & x(705) & x(706) & x(707) & x(708) & x(709) & x(711) & x(712) & x(719) & x(721) & x(725) & x(726) & x(734) & x(735) & x(736) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(750) & x(753) & x(757) & x(761) & x(764) & x(765) & x(766) & x(769) & x(770) & x(771) & x(772) & x(773) & x(774);
    y(23) <= not(p23_out);
    p23 : perceptron
        Generic map (
            WEIGHTS => "111111111100100011111101110111000000000000000001000001000011011000011100111111111111111111111111000001000000000110000000000110000000000",
            SHIFT => 4,
            B => 142,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p23_in,
            y(0) => p23_out,
            y(1 to 17 - 1) => dummy23
        );


    p24_in <= x(40) & x(78) & x(105) & x(126) & x(127) & x(210) & x(238) & x(248) & x(259) & x(260) & x(266) & x(287) & x(289) & x(294) & x(295) & x(320) & x(330) & x(339) & x(346) & x(347) & x(348) & x(349) & x(360) & x(361) & x(366) & x(375) & x(376) & x(377) & x(388) & x(450) & x(474) & x(501) & x(502) & x(509) & x(526) & x(529) & x(534) & x(538) & x(553) & x(584) & x(638) & x(656) & x(657) & x(658) & x(666) & x(675) & x(737) & x(738) & x(739) & x(742) & x(746) & x(747) & x(764);
    y(24) <= not(p24_out);
    p24 : perceptron
        Generic map (
            WEIGHTS => "11100001110110011011111101111100000010000111010000000",
            SHIFT => 4,
            B => -136,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p24_in,
            y(0) => p24_out,
            y(1 to 15 - 1) => dummy24
        );


    p25_in <= x(73) & x(165) & x(166) & x(185) & x(192) & x(193) & x(198) & x(220) & x(221) & x(244) & x(247) & x(248) & x(249) & x(250) & x(266) & x(276) & x(277) & x(278) & x(293) & x(294) & x(295) & x(304) & x(305) & x(306) & x(307) & x(309) & x(320) & x(334) & x(338) & x(339) & x(346) & x(347) & x(348) & x(349) & x(361) & x(366) & x(374) & x(375) & x(376) & x(416) & x(444) & x(450) & x(469) & x(473) & x(474) & x(478) & x(489) & x(490) & x(495) & x(497) & x(501) & x(502) & x(506) & x(516) & x(517) & x(528) & x(529) & x(530) & x(534) & x(545) & x(550) & x(556) & x(557) & x(558) & x(577) & x(584) & x(611) & x(612) & x(638) & x(640) & x(647) & x(648) & x(649) & x(656) & x(657) & x(674) & x(675) & x(676) & x(677) & x(678) & x(712) & x(716) & x(717) & x(718) & x(740) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(770) & x(773);
    y(25) <= not(p25_out);
    p25 : perceptron
        Generic map (
            WEIGHTS => "111111011111110111000111101100111110111111100100110010000010100010000011111111110000000000000",
            SHIFT => 4,
            B => 83,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p25_in,
            y(0) => p25_out,
            y(1 to 16 - 1) => dummy25
        );


    p26_in <= x(63) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(92) & x(95) & x(97) & x(98) & x(99) & x(123) & x(124) & x(125) & x(126) & x(127) & x(162) & x(163) & x(182) & x(183) & x(184) & x(190) & x(191) & x(200) & x(209) & x(210) & x(211) & x(212) & x(219) & x(221) & x(228) & x(238) & x(248) & x(249) & x(250) & x(276) & x(277) & x(278) & x(297) & x(305) & x(306) & x(309) & x(311) & x(333) & x(422) & x(450) & x(509) & x(526) & x(557) & x(692) & x(693) & x(694) & x(695) & x(709) & x(710) & x(711) & x(712) & x(713) & x(715) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(739) & x(742) & x(744) & x(745) & x(746) & x(747) & x(748) & x(749);
    y(26) <= not(p26_out);
    p26 : perceptron
        Generic map (
            WEIGHTS => "1111111111111111100111000111101011111110110010011011111111111111111111111111",
            SHIFT => 4,
            B => 899,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p26_in,
            y(0) => p26_out,
            y(1 to 16 - 1) => dummy26
        );


    p27_in <= x(35) & x(36) & x(37) & x(38) & x(39) & x(40) & x(41) & x(44) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(78) & x(79) & x(90) & x(91) & x(92) & x(93) & x(94) & x(95) & x(96) & x(97) & x(98) & x(99) & x(100) & x(101) & x(102) & x(103) & x(104) & x(105) & x(106) & x(124) & x(135) & x(136) & x(162) & x(163) & x(164) & x(191) & x(192) & x(193) & x(219) & x(220) & x(248) & x(263) & x(277) & x(341) & x(342) & x(368) & x(369) & x(370) & x(371) & x(396) & x(397) & x(398) & x(417) & x(425) & x(445) & x(473) & x(474) & x(479) & x(501) & x(502) & x(507) & x(514) & x(515) & x(529) & x(541) & x(542) & x(543) & x(544) & x(557) & x(563) & x(564) & x(570) & x(591) & x(592) & x(619) & x(620) & x(647) & x(693) & x(694) & x(708) & x(773);
    y(27) <= not(p27_out);
    p27 : perceptron
        Generic map (
            WEIGHTS => "1111111111111111111111111111111111111111111000000000000000000000010111111111111111111111110000",
            SHIFT => 4,
            B => 669,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p27_in,
            y(0) => p27_out,
            y(1 to 16 - 1) => dummy27
        );


    p28_in <= x(35) & x(36) & x(37) & x(38) & x(39) & x(40) & x(41) & x(42) & x(44) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(77) & x(78) & x(79) & x(90) & x(91) & x(92) & x(93) & x(94) & x(95) & x(96) & x(97) & x(103) & x(104) & x(105) & x(106) & x(171) & x(182) & x(197) & x(199) & x(210) & x(211) & x(238) & x(249) & x(276) & x(277) & x(297) & x(299) & x(302) & x(307) & x(332) & x(333) & x(360) & x(361) & x(397) & x(422) & x(424) & x(425) & x(445) & x(450) & x(473) & x(474) & x(501) & x(502) & x(515) & x(529) & x(542) & x(543) & x(557) & x(584) & x(638) & x(640) & x(666) & x(675) & x(694) & x(709) & x(710) & x(712) & x(713) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(732) & x(738) & x(739) & x(740) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(748) & x(749) & x(773);
    y(28) <= not(p28_out);
    p28 : perceptron
        Generic map (
            WEIGHTS => "1111111111111111111111111111111111111101001111110000000000001011111111111110111111111111111111111111110",
            SHIFT => 5,
            B => 1898,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p28_in,
            y(0) => p28_out,
            y(1 to 17 - 1) => dummy28
        );


    p29_in <= x(66) & x(146) & x(155) & x(210) & x(211) & x(221) & x(222) & x(248) & x(249) & x(250) & x(276) & x(277) & x(278) & x(289) & x(330) & x(331) & x(332) & x(341) & x(342) & x(358) & x(359) & x(360) & x(366) & x(387) & x(388) & x(433) & x(453) & x(454) & x(513) & x(514) & x(515) & x(590) & x(591) & x(619) & x(677) & x(692) & x(694) & x(706) & x(707) & x(708) & x(709) & x(710) & x(711) & x(712) & x(715) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(739) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(748) & x(764) & x(770) & x(773);
    y(29) <= not(p29_out);
    p29 : perceptron
        Generic map (
            WEIGHTS => "0110000000000011100111011111111111000000000000000000000000000000",
            SHIFT => 5,
            B => -697,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p29_in,
            y(0) => p29_out,
            y(1 to 17 - 1) => dummy29
        );


    p30_in <= x(41) & x(68) & x(70) & x(74) & x(75) & x(76) & x(77) & x(78) & x(79) & x(100) & x(101) & x(102) & x(103) & x(104) & x(105) & x(106) & x(107) & x(108) & x(138) & x(165) & x(166) & x(182) & x(192) & x(193) & x(194) & x(198) & x(220) & x(221) & x(222) & x(227) & x(244) & x(245) & x(246) & x(247) & x(248) & x(249) & x(250) & x(251) & x(275) & x(276) & x(277) & x(278) & x(289) & x(295) & x(297) & x(298) & x(304) & x(305) & x(306) & x(307) & x(309) & x(310) & x(311) & x(315) & x(333) & x(334) & x(337) & x(338) & x(339) & x(347) & x(348) & x(349) & x(350) & x(361) & x(362) & x(366) & x(376) & x(377) & x(378) & x(386) & x(387) & x(389) & x(390) & x(391) & x(406) & x(418) & x(433) & x(461) & x(501) & x(517) & x(529) & x(544) & x(545) & x(546) & x(557) & x(584) & x(655) & x(656) & x(657) & x(659) & x(681) & x(682) & x(685) & x(692) & x(694) & x(695) & x(706) & x(707) & x(708) & x(719) & x(720) & x(721) & x(722) & x(723) & x(735) & x(736) & x(738) & x(739) & x(741) & x(742) & x(743) & x(748) & x(749) & x(764) & x(765) & x(769) & x(770) & x(771) & x(772) & x(773) & x(774);
    y(30) <= not(p30_out);
    p30 : perceptron
        Generic map (
            WEIGHTS => "1111111111111111110000000100010000000000000111000011100011100000010001100000001111111100000000001110000011111110011111111",
            SHIFT => 4,
            B => 62,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p30_in,
            y(0) => p30_out,
            y(1 to 17 - 1) => dummy30
        );


    p31_in <= x(63) & x(64) & x(91) & x(92) & x(93) & x(98) & x(99) & x(106) & x(108) & x(147) & x(151) & x(165) & x(166) & x(171) & x(172) & x(175) & x(176) & x(177) & x(178) & x(179) & x(180) & x(192) & x(193) & x(199) & x(200) & x(201) & x(210) & x(211) & x(213) & x(220) & x(221) & x(222) & x(247) & x(248) & x(249) & x(250) & x(276) & x(277) & x(296) & x(297) & x(298) & x(299) & x(300) & x(301) & x(302) & x(305) & x(306) & x(309) & x(324) & x(325) & x(327) & x(328) & x(330) & x(331) & x(332) & x(334) & x(350) & x(359) & x(360) & x(388) & x(406) & x(416) & x(433) & x(436) & x(450) & x(455) & x(456) & x(461) & x(488) & x(489) & x(490) & x(493) & x(506) & x(517) & x(518) & x(534) & x(535) & x(583) & x(611) & x(619) & x(647) & x(648) & x(655) & x(675) & x(676) & x(677) & x(678) & x(679) & x(706) & x(708) & x(719) & x(720) & x(721) & x(746) & x(747) & x(748);
    y(31) <= not(p31_out);
    p31 : perceptron
        Generic map (
            WEIGHTS => "000001111110011111111001111110000000001111111001111111100111010111100001100110011111111111111111",
            SHIFT => 4,
            B => 327,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p31_in,
            y(0) => p31_out,
            y(1 to 16 - 1) => dummy31
        );


    p32_in <= x(37) & x(45) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(90) & x(91) & x(92) & x(210) & x(211) & x(221) & x(222) & x(238) & x(248) & x(249) & x(250) & x(276) & x(277) & x(278) & x(299) & x(300) & x(301) & x(302) & x(303) & x(304) & x(305) & x(311) & x(327) & x(329) & x(330) & x(331) & x(332) & x(340) & x(358) & x(359) & x(360) & x(361) & x(368) & x(424) & x(425) & x(453) & x(485) & x(513) & x(514) & x(534) & x(657) & x(658) & x(677) & x(694) & x(709) & x(710) & x(711) & x(712) & x(713) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(737) & x(738) & x(739) & x(740) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(748) & x(749);
    y(32) <= not(p32_out);
    p32 : perceptron
        Generic map (
            WEIGHTS => "00000000000000000000000011111101111110111101111111110000000000000000000000000000",
            SHIFT => 4,
            B => -730,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p32_in,
            y(0) => p32_out,
            y(1 to 16 - 1) => dummy32
        );


    p33_in <= x(0) & x(1) & x(2) & x(3) & x(4) & x(5) & x(6) & x(7) & x(8) & x(9) & x(10) & x(11) & x(12) & x(15) & x(16) & x(17) & x(18) & x(19) & x(20) & x(21) & x(22) & x(23) & x(24) & x(25) & x(26) & x(27) & x(28) & x(29) & x(30) & x(31) & x(35) & x(39) & x(40) & x(41) & x(43) & x(52) & x(53) & x(54) & x(55) & x(56) & x(57) & x(58) & x(59) & x(63) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(79) & x(82) & x(83) & x(84) & x(85) & x(87) & x(88) & x(96) & x(97) & x(98) & x(99) & x(101) & x(102) & x(103) & x(104) & x(105) & x(106) & x(107) & x(108) & x(110) & x(111) & x(112) & x(115) & x(139) & x(141) & x(142) & x(167) & x(169) & x(193) & x(196) & x(197) & x(200) & x(238) & x(239) & x(248) & x(260) & x(261) & x(266) & x(267) & x(275) & x(276) & x(294) & x(295) & x(303) & x(304) & x(320) & x(322) & x(323) & x(330) & x(331) & x(332) & x(345) & x(347) & x(348) & x(349) & x(353) & x(359) & x(360) & x(364) & x(375) & x(376) & x(380) & x(381) & x(388) & x(389) & x(392) & x(403) & x(408) & x(416) & x(419) & x(420) & x(432) & x(436) & x(444) & x(449) & x(450) & x(463) & x(476) & x(478) & x(489) & x(501) & x(502) & x(503) & x(504) & x(506) & x(517) & x(528) & x(529) & x(530) & x(532) & x(534) & x(556) & x(557) & x(558) & x(560) & x(583) & x(584) & x(585) & x(587) & x(588) & x(611) & x(612) & x(615) & x(616) & x(617) & x(618) & x(638) & x(639) & x(643) & x(644) & x(645) & x(647) & x(656) & x(671) & x(672) & x(673) & x(675) & x(679) & x(692) & x(693) & x(695) & x(699) & x(700) & x(701) & x(702) & x(709) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(724) & x(725) & x(726) & x(727) & x(728) & x(729) & x(730) & x(731) & x(747) & x(748) & x(749) & x(752) & x(753) & x(755) & x(756) & x(757) & x(758) & x(759) & x(760) & x(779) & x(781) & x(782) & x(783);
    y(33) <= not(p33_out);
    p33 : perceptron
        Generic map (
            WEIGHTS => "000000000000000000000000000000111110000000011111111111111100000011111111111100000000010110011100110011100111111111101111110111001110110100000100000100000000000000100000110001111100001111111110000000111000000000000",
            SHIFT => 4,
            B => -648,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p33_in,
            y(0) => p33_out,
            y(1 to 17 - 1) => dummy33
        );


    p34_in <= x(2) & x(11) & x(15) & x(30) & x(53) & x(56) & x(58) & x(63) & x(64) & x(67) & x(68) & x(70) & x(75) & x(76) & x(78) & x(79) & x(91) & x(93) & x(94) & x(95) & x(96) & x(97) & x(98) & x(99) & x(100) & x(101) & x(102) & x(103) & x(104) & x(105) & x(106) & x(107) & x(108) & x(140) & x(165) & x(166) & x(191) & x(192) & x(193) & x(194) & x(196) & x(219) & x(220) & x(221) & x(222) & x(247) & x(248) & x(249) & x(250) & x(276) & x(277) & x(278) & x(289) & x(294) & x(295) & x(298) & x(305) & x(306) & x(307) & x(309) & x(310) & x(316) & x(317) & x(319) & x(321) & x(328) & x(329) & x(330) & x(333) & x(334) & x(337) & x(338) & x(346) & x(347) & x(348) & x(349) & x(350) & x(357) & x(358) & x(361) & x(362) & x(366) & x(375) & x(376) & x(377) & x(378) & x(381) & x(394) & x(406) & x(408) & x(409) & x(419) & x(449) & x(465) & x(473) & x(474) & x(501) & x(502) & x(514) & x(515) & x(517) & x(529) & x(544) & x(545) & x(557) & x(584) & x(612) & x(644) & x(646) & x(655) & x(656) & x(657) & x(660) & x(671) & x(682) & x(684) & x(699) & x(703) & x(706) & x(707) & x(708) & x(709) & x(716) & x(717) & x(718) & x(719) & x(721) & x(732) & x(735) & x(736) & x(737) & x(738) & x(739) & x(740) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(748) & x(755) & x(769) & x(770) & x(772) & x(773) & x(774) & x(775);
    y(34) <= not(p34_out);
    p34 : perceptron
        Generic map (
            WEIGHTS => "11111110000000000000000000000000011111111111111111111000111001111000110011111001101111101111110000000000000111111111110000000000000000000000001000000",
            SHIFT => 4,
            B => -362,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p34_in,
            y(0) => p34_out,
            y(1 to 17 - 1) => dummy34
        );


    p35_in <= x(0) & x(1) & x(2) & x(3) & x(4) & x(5) & x(6) & x(7) & x(8) & x(9) & x(10) & x(11) & x(12) & x(15) & x(16) & x(17) & x(18) & x(19) & x(20) & x(21) & x(22) & x(23) & x(24) & x(25) & x(26) & x(27) & x(28) & x(29) & x(30) & x(31) & x(32) & x(33) & x(35) & x(37) & x(39) & x(40) & x(44) & x(52) & x(53) & x(54) & x(55) & x(56) & x(57) & x(58) & x(59) & x(61) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(79) & x(82) & x(83) & x(84) & x(85) & x(87) & x(88) & x(90) & x(91) & x(92) & x(93) & x(94) & x(95) & x(96) & x(97) & x(98) & x(100) & x(105) & x(110) & x(111) & x(112) & x(113) & x(115) & x(121) & x(122) & x(138) & x(139) & x(140) & x(141) & x(142) & x(167) & x(168) & x(169) & x(196) & x(221) & x(222) & x(248) & x(249) & x(250) & x(276) & x(277) & x(278) & x(297) & x(298) & x(299) & x(300) & x(301) & x(302) & x(303) & x(305) & x(306) & x(329) & x(330) & x(331) & x(332) & x(340) & x(359) & x(360) & x(364) & x(367) & x(387) & x(388) & x(392) & x(397) & x(416) & x(417) & x(419) & x(420) & x(424) & x(425) & x(445) & x(448) & x(449) & x(451) & x(453) & x(473) & x(474) & x(476) & x(479) & x(501) & x(503) & x(504) & x(507) & x(529) & x(532) & x(535) & x(560) & x(563) & x(587) & x(588) & x(615) & x(616) & x(617) & x(643) & x(644) & x(645) & x(671) & x(672) & x(673) & x(698) & x(699) & x(700) & x(701) & x(702) & x(708) & x(709) & x(710) & x(711) & x(712) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(725) & x(726) & x(727) & x(728) & x(729) & x(730) & x(731) & x(734) & x(737) & x(738) & x(739) & x(740) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(748) & x(749) & x(750) & x(752) & x(753) & x(754) & x(755) & x(756) & x(757) & x(758) & x(759) & x(760) & x(770) & x(779) & x(780) & x(781) & x(782) & x(783);
    y(35) <= not(p35_out);
    p35 : perceptron
        Generic map (
            WEIGHTS => "11111111111111111111111111111111000001111111110000000000011111100000000000111110001111111100000000111111100111101110111110111101101001001100101011111111111111110000000000001111111000000000000000111111111011111",
            SHIFT => 5,
            B => 1022,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p35_in,
            y(0) => p35_out,
            y(1 to 18 - 1) => dummy35
        );


    p36_in <= x(39) & x(40) & x(41) & x(42) & x(43) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(102) & x(103) & x(104) & x(105) & x(106) & x(107) & x(108) & x(162) & x(171) & x(172) & x(248) & x(255) & x(264) & x(265) & x(269) & x(276) & x(283) & x(284) & x(292) & x(295) & x(304) & x(320) & x(321) & x(322) & x(339) & x(347) & x(348) & x(349) & x(350) & x(351) & x(352) & x(376) & x(377) & x(388) & x(389) & x(406) & x(407) & x(416) & x(433) & x(434) & x(446) & x(450) & x(460) & x(462) & x(473) & x(474) & x(501) & x(502) & x(506) & x(509) & x(510) & x(511) & x(518) & x(528) & x(529) & x(530) & x(534) & x(535) & x(539) & x(545) & x(556) & x(557) & x(558) & x(562) & x(583) & x(584) & x(611) & x(612) & x(637) & x(638) & x(639) & x(640) & x(647) & x(656) & x(657) & x(675) & x(682) & x(693) & x(695) & x(709) & x(711) & x(712) & x(713) & x(719) & x(720) & x(721) & x(722) & x(723) & x(724) & x(735) & x(736) & x(740) & x(742) & x(748) & x(749) & x(769) & x(771) & x(772);
    y(36) <= not(p36_out);
    p36 : perceptron
        Generic map (
            WEIGHTS => "11111111111111111111111110111000010000111101111111111111110111000010000000110000010000000011111110000111111000011000",
            SHIFT => 4,
            B => 260,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p36_in,
            y(0) => p36_out,
            y(1 to 16 - 1) => dummy36
        );


    p37_in <= x(40) & x(43) & x(65) & x(66) & x(67) & x(68) & x(69) & x(71) & x(73) & x(137) & x(138) & x(165) & x(166) & x(188) & x(192) & x(193) & x(194) & x(198) & x(220) & x(221) & x(222) & x(226) & x(248) & x(249) & x(250) & x(251) & x(276) & x(277) & x(278) & x(296) & x(297) & x(298) & x(299) & x(300) & x(305) & x(306) & x(309) & x(310) & x(311) & x(322) & x(324) & x(326) & x(328) & x(329) & x(333) & x(334) & x(337) & x(338) & x(339) & x(348) & x(349) & x(350) & x(351) & x(355) & x(356) & x(366) & x(376) & x(377) & x(378) & x(406) & x(433) & x(450) & x(451) & x(461) & x(478) & x(479) & x(486) & x(501) & x(502) & x(506) & x(507) & x(513) & x(514) & x(528) & x(529) & x(530) & x(534) & x(535) & x(556) & x(557) & x(558) & x(563) & x(584) & x(591) & x(612) & x(619) & x(625) & x(638) & x(646) & x(647) & x(648) & x(654) & x(674) & x(675) & x(676) & x(677) & x(678) & x(693) & x(694) & x(695) & x(704) & x(719) & x(720) & x(721) & x(722) & x(723) & x(724) & x(735) & x(748) & x(749) & x(769) & x(770) & x(773) & x(774);
    y(37) <= not(p37_out);
    p37 : perceptron
        Generic map (
            WEIGHTS => "000000000000000001000100000001111100111011110011100001110000000000111001111100111010100100000000000010000001001111",
            SHIFT => 4,
            B => -536,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p37_in,
            y(0) => p37_out,
            y(1 to 16 - 1) => dummy37
        );


    p38_in <= x(37) & x(40) & x(135) & x(188) & x(192) & x(221) & x(222) & x(227) & x(248) & x(249) & x(250) & x(277) & x(302) & x(303) & x(322) & x(323) & x(326) & x(328) & x(329) & x(330) & x(331) & x(332) & x(342) & x(350) & x(357) & x(358) & x(359) & x(360) & x(368) & x(369) & x(370) & x(378) & x(390) & x(418) & x(429) & x(446) & x(450) & x(453) & x(454) & x(473) & x(474) & x(481) & x(485) & x(486) & x(501) & x(502) & x(512) & x(513) & x(514) & x(515) & x(528) & x(529) & x(535) & x(542) & x(547) & x(556) & x(557) & x(558) & x(584) & x(612) & x(640) & x(648) & x(652) & x(653) & x(675) & x(676) & x(677) & x(678) & x(679) & x(694) & x(705) & x(706) & x(707) & x(708) & x(709);
    y(38) <= not(p38_out);
    p38 : perceptron
        Generic map (
            WEIGHTS => "000000000000110011111100111100001111011111111111111101111111100000000000000",
            SHIFT => 4,
            B => 8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p38_in,
            y(0) => p38_out,
            y(1 to 16 - 1) => dummy38
        );


    p39_in <= x(44) & x(64) & x(66) & x(67) & x(68) & x(69) & x(70) & x(75) & x(76) & x(91) & x(93) & x(94) & x(95) & x(96) & x(100) & x(101) & x(102) & x(103) & x(104) & x(108) & x(136) & x(171) & x(172) & x(210) & x(211) & x(213) & x(249) & x(304) & x(311) & x(332) & x(333) & x(339) & x(341) & x(342) & x(349) & x(350) & x(369) & x(377) & x(379) & x(380) & x(406) & x(407) & x(414) & x(433) & x(445) & x(450) & x(461) & x(468) & x(473) & x(482) & x(500) & x(501) & x(502) & x(506) & x(511) & x(528) & x(529) & x(530) & x(534) & x(544) & x(545) & x(549) & x(555) & x(556) & x(557) & x(558) & x(575) & x(576) & x(583) & x(584) & x(602) & x(610) & x(611) & x(612) & x(637) & x(638) & x(639) & x(640) & x(647) & x(675) & x(676) & x(677) & x(692) & x(693) & x(694) & x(695) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(724) & x(745) & x(746) & x(747) & x(748) & x(749);
    y(39) <= not(p39_out);
    p39 : perceptron
        Generic map (
            WEIGHTS => "0000000000000000000111111111011011111111110101100000010000100000000000000000001111111111111111111111",
            SHIFT => 4,
            B => -88,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p39_in,
            y(0) => p39_out,
            y(1 to 16 - 1) => dummy39
        );


    p40_in <= x(35) & x(37) & x(38) & x(39) & x(40) & x(44) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(78) & x(79) & x(90) & x(91) & x(92) & x(93) & x(94) & x(95) & x(96) & x(97) & x(104) & x(105) & x(154) & x(156) & x(157) & x(181) & x(184) & x(198) & x(199) & x(206) & x(219) & x(220) & x(221) & x(227) & x(247) & x(248) & x(249) & x(276) & x(277) & x(295) & x(297) & x(299) & x(322) & x(323) & x(325) & x(327) & x(348) & x(350) & x(361) & x(366) & x(376) & x(403) & x(411) & x(418) & x(423) & x(437) & x(459) & x(501) & x(526) & x(527) & x(529) & x(539) & x(541) & x(542) & x(543) & x(549) & x(557) & x(566) & x(569) & x(581) & x(582) & x(584) & x(595) & x(599) & x(606) & x(611) & x(707) & x(718) & x(735) & x(736) & x(737) & x(744) & x(746) & x(773);
    y(40) <= not(p40_out);
    p40 : perceptron
        Generic map (
            WEIGHTS => "11111111111111111111111111111111001111011111000000010001100001111111111111111111100000000",
            SHIFT => 4,
            B => 479,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p40_in,
            y(0) => p40_out,
            y(1 to 16 - 1) => dummy40
        );


    p41_in <= x(62) & x(63) & x(64) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(90) & x(91) & x(92) & x(93) & x(98) & x(101) & x(102) & x(103) & x(104) & x(106) & x(107) & x(108) & x(166) & x(171) & x(172) & x(173) & x(174) & x(187) & x(193) & x(199) & x(200) & x(220) & x(221) & x(227) & x(228) & x(247) & x(248) & x(249) & x(250) & x(275) & x(276) & x(277) & x(295) & x(297) & x(298) & x(299) & x(300) & x(306) & x(309) & x(324) & x(326) & x(360) & x(385) & x(416) & x(433) & x(441) & x(450) & x(460) & x(501) & x(506) & x(534) & x(535) & x(542) & x(563) & x(569) & x(583) & x(598) & x(610) & x(611) & x(619) & x(638) & x(640) & x(647) & x(648) & x(675) & x(676) & x(677) & x(678) & x(679) & x(705) & x(706) & x(707) & x(708) & x(736) & x(743) & x(770) & x(773);
    y(41) <= not(p41_out);
    p41 : perceptron
        Generic map (
            WEIGHTS => "000111111100001111111101111001100110000000111110111111011001110100000100111111111111111",
            SHIFT => 5,
            B => 580,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p41_in,
            y(0) => p41_out,
            y(1 to 17 - 1) => dummy41
        );


    p42_in <= x(37) & x(45) & x(46) & x(49) & x(64) & x(68) & x(70) & x(73) & x(75) & x(78) & x(79) & x(104) & x(105) & x(108) & x(135) & x(163) & x(164) & x(165) & x(183) & x(191) & x(192) & x(193) & x(194) & x(197) & x(210) & x(211) & x(219) & x(220) & x(221) & x(222) & x(238) & x(248) & x(249) & x(250) & x(276) & x(277) & x(278) & x(279) & x(283) & x(301) & x(302) & x(303) & x(304) & x(305) & x(312) & x(326) & x(328) & x(329) & x(330) & x(331) & x(332) & x(347) & x(350) & x(355) & x(356) & x(357) & x(358) & x(359) & x(360) & x(400) & x(418) & x(422) & x(446) & x(450) & x(472) & x(479) & x(484) & x(485) & x(487) & x(507) & x(513) & x(514) & x(515) & x(516) & x(534) & x(535) & x(542) & x(543) & x(563) & x(584) & x(591) & x(618) & x(619) & x(647) & x(648) & x(675) & x(676) & x(677) & x(678) & x(690) & x(691) & x(692) & x(693) & x(695) & x(703) & x(704) & x(705) & x(706) & x(707) & x(708) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(735) & x(745) & x(746) & x(747) & x(748) & x(749) & x(765) & x(766) & x(767) & x(768) & x(769) & x(770) & x(771) & x(773);
    y(42) <= not(p42_out);
    p42 : perceptron
        Generic map (
            WEIGHTS => "11111111111110111101111100111101111111100001100000010000000101011100010000110011111111111000001111110000000010000011111111",
            SHIFT => 4,
            B => 566,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p42_in,
            y(0) => p42_out,
            y(1 to 17 - 1) => dummy42
        );


    p43_in <= x(96) & x(105) & x(123) & x(124) & x(125) & x(126) & x(127) & x(151) & x(152) & x(153) & x(162) & x(163) & x(181) & x(182) & x(183) & x(184) & x(185) & x(189) & x(190) & x(191) & x(198) & x(210) & x(211) & x(212) & x(213) & x(219) & x(226) & x(238) & x(239) & x(240) & x(248) & x(249) & x(250) & x(254) & x(276) & x(277) & x(278) & x(282) & x(284) & x(288) & x(291) & x(293) & x(304) & x(306) & x(309) & x(310) & x(311) & x(312) & x(316) & x(318) & x(338) & x(339) & x(343) & x(344) & x(346) & x(347) & x(350) & x(366) & x(371) & x(374) & x(378) & x(390) & x(391) & x(450) & x(479) & x(507) & x(534) & x(535) & x(563) & x(564) & x(591) & x(619) & x(620) & x(647) & x(648) & x(674) & x(675) & x(693) & x(694) & x(695) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(732) & x(746) & x(747) & x(748) & x(749) & x(764) & x(765) & x(769) & x(770) & x(771) & x(772) & x(773) & x(774);
    y(43) <= not(p43_out);
    p43 : perceptron
        Generic map (
            WEIGHTS => "01000000001100000111100001100000010001111100111111111111011100000000000000000000000000000000011111111",
            SHIFT => 4,
            B => -236,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p43_in,
            y(0) => p43_out,
            y(1 to 16 - 1) => dummy43
        );


    p44_in <= x(37) & x(38) & x(39) & x(40) & x(41) & x(45) & x(46) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(79) & x(101) & x(102) & x(103) & x(104) & x(105) & x(106) & x(107) & x(108) & x(147) & x(158) & x(171) & x(172) & x(186) & x(187) & x(188) & x(238) & x(246) & x(249) & x(266) & x(305) & x(352) & x(362) & x(375) & x(381) & x(390) & x(399) & x(400) & x(408) & x(409) & x(411) & x(414) & x(418) & x(423) & x(436) & x(437) & x(446) & x(450) & x(451) & x(464) & x(473) & x(474) & x(478) & x(481) & x(501) & x(502) & x(506) & x(507) & x(528) & x(529) & x(534) & x(535) & x(557) & x(562) & x(563) & x(576) & x(584) & x(591) & x(597) & x(598) & x(618) & x(619) & x(638) & x(647) & x(648) & x(649) & x(659) & x(675) & x(676) & x(677) & x(678) & x(679) & x(705) & x(706) & x(708);
    y(44) <= not(p44_out);
    p44 : perceptron
        Generic map (
            WEIGHTS => "11111111111111111111111111111111101100000001101101111110111011100100011001101110100110111011111111",
            SHIFT => 4,
            B => 846,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p44_in,
            y(0) => p44_out,
            y(1 to 16 - 1) => dummy44
        );


    p45_in <= x(73) & x(76) & x(78) & x(104) & x(105) & x(106) & x(149) & x(150) & x(160) & x(198) & x(199) & x(226) & x(227) & x(228) & x(249) & x(250) & x(254) & x(255) & x(256) & x(266) & x(267) & x(268) & x(269) & x(270) & x(281) & x(282) & x(283) & x(284) & x(294) & x(295) & x(309) & x(310) & x(311) & x(312) & x(338) & x(339) & x(348) & x(353) & x(358) & x(359) & x(360) & x(361) & x(362) & x(366) & x(367) & x(376) & x(377) & x(378) & x(380) & x(390) & x(403) & x(404) & x(405) & x(415) & x(418) & x(424) & x(431) & x(432) & x(433) & x(436) & x(446) & x(460) & x(474) & x(482) & x(483) & x(487) & x(488) & x(514) & x(515) & x(535) & x(571) & x(676) & x(677) & x(678) & x(692) & x(693) & x(694) & x(695) & x(696) & x(706) & x(707) & x(708) & x(718) & x(719) & x(720) & x(721) & x(722) & x(732) & x(735) & x(736) & x(737) & x(743) & x(748) & x(749) & x(764) & x(765) & x(766) & x(768) & x(769) & x(770) & x(771) & x(772) & x(773) & x(774);
    y(45) <= not(p45_out);
    p45 : perceptron
        Generic map (
            WEIGHTS => "00000000111111111111111111111111111100000111100001000110000010111000011111000001110000001111001111111111",
            SHIFT => 4,
            B => 314,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p45_in,
            y(0) => p45_out,
            y(1 to 16 - 1) => dummy45
        );


    p46_in <= x(35) & x(39) & x(63) & x(64) & x(66) & x(67) & x(68) & x(70) & x(79) & x(94) & x(126) & x(127) & x(135) & x(136) & x(164) & x(171) & x(172) & x(192) & x(198) & x(199) & x(200) & x(201) & x(202) & x(210) & x(211) & x(212) & x(218) & x(227) & x(228) & x(229) & x(238) & x(239) & x(249) & x(254) & x(255) & x(256) & x(259) & x(270) & x(283) & x(284) & x(294) & x(295) & x(298) & x(305) & x(307) & x(310) & x(312) & x(322) & x(323) & x(324) & x(326) & x(333) & x(334) & x(339) & x(350) & x(351) & x(358) & x(359) & x(360) & x(361) & x(362) & x(366) & x(387) & x(388) & x(394) & x(402) & x(403) & x(422) & x(423) & x(429) & x(430) & x(431) & x(434) & x(435) & x(438) & x(450) & x(451) & x(458) & x(461) & x(462) & x(483) & x(486) & x(501) & x(502) & x(507) & x(513) & x(514) & x(528) & x(529) & x(535) & x(538) & x(542) & x(543) & x(552) & x(554) & x(556) & x(557) & x(568) & x(576) & x(584) & x(612) & x(638) & x(666) & x(677) & x(678) & x(679) & x(697) & x(706) & x(707) & x(708) & x(721) & x(735) & x(736) & x(737) & x(742) & x(743) & x(744) & x(748) & x(764) & x(765) & x(769) & x(770) & x(773) & x(774);
    y(46) <= not(p46_out);
    p46 : perceptron
        Generic map (
            WEIGHTS => "1111111111110000000000011100001100000000000000000000000011100011011001110000010011110111101111111111111000100010000001000000",
            SHIFT => 4,
            B => -301,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p46_in,
            y(0) => p46_out,
            y(1 to 17 - 1) => dummy46
        );


    p47_in <= x(63) & x(64) & x(124) & x(151) & x(153) & x(154) & x(165) & x(166) & x(190) & x(191) & x(192) & x(193) & x(198) & x(210) & x(219) & x(220) & x(221) & x(226) & x(238) & x(247) & x(248) & x(249) & x(250) & x(262) & x(276) & x(277) & x(288) & x(289) & x(291) & x(295) & x(315) & x(319) & x(320) & x(323) & x(332) & x(345) & x(347) & x(348) & x(350) & x(372) & x(373) & x(390) & x(473) & x(474) & x(479) & x(502) & x(507) & x(529) & x(535) & x(557) & x(563) & x(591) & x(618) & x(619) & x(620) & x(623) & x(624) & x(647) & x(648) & x(719) & x(720) & x(721) & x(723) & x(748);
    y(47) <= not(p47_out);
    p47 : perceptron
        Generic map (
            WEIGHTS => "1100001111111011110111111111101110011101100000000000000000000000",
            SHIFT => 4,
            B => -65,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p47_in,
            y(0) => p47_out,
            y(1 to 16 - 1) => dummy47
        );


    p48_in <= x(37) & x(38) & x(39) & x(40) & x(41) & x(43) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(102) & x(103) & x(104) & x(105) & x(106) & x(118) & x(121) & x(123) & x(125) & x(133) & x(150) & x(151) & x(153) & x(180) & x(182) & x(183) & x(184) & x(186) & x(210) & x(211) & x(212) & x(213) & x(240) & x(243) & x(244) & x(259) & x(287) & x(302) & x(303) & x(304) & x(331) & x(332) & x(361) & x(362) & x(386) & x(387) & x(390) & x(391) & x(412) & x(414) & x(418) & x(446) & x(450) & x(453) & x(473) & x(474) & x(479) & x(490) & x(501) & x(502) & x(507) & x(528) & x(529) & x(530) & x(535) & x(539) & x(545) & x(553) & x(554) & x(556) & x(557) & x(558) & x(563) & x(564) & x(565) & x(566) & x(567) & x(568) & x(572) & x(574) & x(584) & x(585) & x(591) & x(592) & x(601) & x(612) & x(613) & x(619) & x(620) & x(622) & x(638) & x(639) & x(640) & x(647) & x(709) & x(710) & x(717) & x(718) & x(719) & x(720) & x(721) & x(723) & x(732) & x(746) & x(747) & x(748) & x(749);
    y(48) <= not(p48_out);
    p48 : perceptron
        Generic map (
            WEIGHTS => "111111111111111111111111111100001000000000000000110000000110011000000010000000010000000000011000010000000000000000000000",
            SHIFT => 4,
            B => -457,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p48_in,
            y(0) => p48_out,
            y(1 to 17 - 1) => dummy48
        );


    p49_in <= x(35) & x(36) & x(37) & x(38) & x(39) & x(40) & x(41) & x(42) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(79) & x(81) & x(90) & x(91) & x(94) & x(95) & x(96) & x(97) & x(98) & x(99) & x(100) & x(101) & x(102) & x(103) & x(104) & x(105) & x(106) & x(107) & x(108) & x(162) & x(163) & x(164) & x(165) & x(190) & x(191) & x(192) & x(193) & x(194) & x(218) & x(219) & x(220) & x(221) & x(222) & x(247) & x(248) & x(249) & x(250) & x(266) & x(276) & x(277) & x(294) & x(333) & x(334) & x(338) & x(366) & x(369) & x(417) & x(445) & x(515) & x(543) & x(655) & x(656) & x(657) & x(659) & x(674) & x(736) & x(737) & x(738) & x(739) & x(741) & x(742) & x(743) & x(746);
    y(49) <= not(p49_out);
    p49 : perceptron
        Generic map (
            WEIGHTS => "1111111111111111111111111101111111111111111100000000000000000010010011011110000011111111",
            SHIFT => 4,
            B => 648,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p49_in,
            y(0) => p49_out,
            y(1 to 16 - 1) => dummy49
        );


    p50_in <= x(78) & x(104) & x(105) & x(106) & x(195) & x(198) & x(199) & x(221) & x(227) & x(248) & x(249) & x(250) & x(266) & x(276) & x(277) & x(278) & x(283) & x(294) & x(305) & x(312) & x(328) & x(329) & x(330) & x(331) & x(338) & x(339) & x(349) & x(357) & x(358) & x(359) & x(360) & x(362) & x(366) & x(376) & x(377) & x(378) & x(379) & x(386) & x(387) & x(390) & x(404) & x(405) & x(418) & x(432) & x(433) & x(446) & x(460) & x(461) & x(473) & x(474) & x(484) & x(485) & x(486) & x(487) & x(488) & x(500) & x(502) & x(513) & x(514) & x(515) & x(516) & x(535) & x(557) & x(584) & x(676) & x(677) & x(690) & x(691) & x(692) & x(693) & x(694) & x(695) & x(706) & x(707) & x(708) & x(710) & x(711) & x(712) & x(719) & x(720) & x(721) & x(722) & x(735) & x(736) & x(737) & x(743) & x(748) & x(764) & x(765) & x(766) & x(769) & x(770) & x(773) & x(774);
    y(50) <= not(p50_out);
    p50 : perceptron
        Generic map (
            WEIGHTS => "1111000000000000000011110011111001111110110110110011111001111000001111110000001111000010000000",
            SHIFT => 4,
            B => -311,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p50_in,
            y(0) => p50_out,
            y(1 to 16 - 1) => dummy50
        );


    p51_in <= x(63) & x(67) & x(68) & x(70) & x(77) & x(78) & x(93) & x(103) & x(104) & x(105) & x(106) & x(107) & x(108) & x(188) & x(192) & x(198) & x(219) & x(221) & x(222) & x(249) & x(250) & x(261) & x(264) & x(277) & x(290) & x(292) & x(303) & x(305) & x(309) & x(310) & x(311) & x(328) & x(329) & x(330) & x(331) & x(332) & x(338) & x(339) & x(350) & x(353) & x(358) & x(366) & x(367) & x(378) & x(390) & x(394) & x(400) & x(445) & x(450) & x(474) & x(507) & x(513) & x(514) & x(515) & x(523) & x(535) & x(563) & x(565) & x(591) & x(647) & x(648) & x(649) & x(675) & x(676) & x(677) & x(678) & x(707) & x(709) & x(710) & x(711) & x(712) & x(713) & x(714) & x(715) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(735) & x(736) & x(737) & x(738) & x(739) & x(740) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(748) & x(750) & x(764) & x(769) & x(770) & x(771) & x(772) & x(773) & x(774) & x(775);
    y(51) <= not(p51_out);
    p51 : perceptron
        Generic map (
            WEIGHTS => "00000000000001101111100100010000000000100001001010100011111111111100000000000000000000000000000000000000",
            SHIFT => 4,
            B => -919,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p51_in,
            y(0) => p51_out,
            y(1 to 16 - 1) => dummy51
        );


    p52_in <= x(35) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(77) & x(78) & x(97) & x(99) & x(102) & x(103) & x(104) & x(105) & x(106) & x(107) & x(108) & x(163) & x(182) & x(183) & x(191) & x(192) & x(195) & x(203) & x(204) & x(210) & x(211) & x(220) & x(221) & x(238) & x(249) & x(277) & x(303) & x(304) & x(328) & x(329) & x(330) & x(331) & x(332) & x(338) & x(357) & x(358) & x(359) & x(360) & x(366) & x(374) & x(394) & x(400) & x(437) & x(439) & x(465) & x(514) & x(515) & x(535) & x(584) & x(695) & x(703) & x(709) & x(714) & x(715) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(736) & x(737) & x(738) & x(739) & x(740) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(748) & x(749) & x(750);
    y(52) <= not(p52_out);
    p52 : perceptron
        Generic map (
            WEIGHTS => "1111111111111111111011000001100100111111111111101000011001011111111111111111111111111",
            SHIFT => 5,
            B => 1057,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p52_in,
            y(0) => p52_out,
            y(1 to 17 - 1) => dummy52
        );


    p53_in <= x(35) & x(44) & x(63) & x(64) & x(65) & x(66) & x(91) & x(92) & x(93) & x(94) & x(134) & x(135) & x(136) & x(171) & x(172) & x(199) & x(200) & x(201) & x(227) & x(231) & x(232) & x(233) & x(234) & x(238) & x(246) & x(248) & x(249) & x(258) & x(261) & x(276) & x(294) & x(295) & x(303) & x(320) & x(322) & x(323) & x(348) & x(399) & x(400) & x(427) & x(428) & x(440) & x(450) & x(456) & x(473) & x(487) & x(501) & x(502) & x(506) & x(514) & x(515) & x(520) & x(529) & x(535) & x(542) & x(557) & x(655) & x(656) & x(676) & x(677) & x(678) & x(682) & x(683) & x(684) & x(685) & x(686) & x(687) & x(706) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(723) & x(732) & x(748) & x(749) & x(764) & x(773);
    y(53) <= not(p53_out);
    p53 : perceptron
        Generic map (
            WEIGHTS => "11111111110000000001111111111100110010000000111101111011110001111110111111111100",
            SHIFT => 4,
            B => 393,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p53_in,
            y(0) => p53_out,
            y(1 to 16 - 1) => dummy53
        );


    p54_in <= x(75) & x(78) & x(102) & x(103) & x(104) & x(105) & x(106) & x(107) & x(165) & x(166) & x(186) & x(192) & x(193) & x(194) & x(198) & x(220) & x(221) & x(222) & x(247) & x(248) & x(249) & x(250) & x(251) & x(275) & x(276) & x(277) & x(278) & x(304) & x(305) & x(306) & x(307) & x(309) & x(324) & x(326) & x(333) & x(334) & x(348) & x(349) & x(350) & x(361) & x(362) & x(383) & x(390) & x(394) & x(409) & x(411) & x(436) & x(446) & x(457) & x(458) & x(479) & x(491) & x(507) & x(537) & x(541) & x(565) & x(574) & x(627) & x(652) & x(656) & x(657) & x(658) & x(659) & x(660) & x(674) & x(703) & x(706) & x(707) & x(708) & x(716) & x(735) & x(736) & x(737) & x(738) & x(739) & x(740) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(770) & x(772) & x(773);
    y(54) <= not(p54_out);
    p54 : perceptron
        Generic map (
            WEIGHTS => "0000000011111101111111111111111000111111101000010010111101111111110000000000000000000",
            SHIFT => 4,
            B => 118,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p54_in,
            y(0) => p54_out,
            y(1 to 16 - 1) => dummy54
        );


    p55_in <= x(97) & x(98) & x(101) & x(105) & x(164) & x(165) & x(189) & x(190) & x(191) & x(192) & x(193) & x(194) & x(217) & x(219) & x(220) & x(221) & x(222) & x(237) & x(238) & x(239) & x(245) & x(247) & x(248) & x(249) & x(250) & x(266) & x(267) & x(273) & x(276) & x(277) & x(278) & x(295) & x(301) & x(302) & x(303) & x(305) & x(320) & x(328) & x(329) & x(330) & x(331) & x(332) & x(347) & x(348) & x(354) & x(371) & x(375) & x(376) & x(390) & x(398) & x(399) & x(400) & x(418) & x(426) & x(431) & x(432) & x(446) & x(474) & x(502) & x(633) & x(634) & x(712) & x(717) & x(718) & x(719) & x(721) & x(742);
    y(55) <= not(p55_out);
    p55 : perceptron
        Generic map (
            WEIGHTS => "1110000000000000011100000110000111100111110010001000100011100111111",
            SHIFT => 4,
            B => -181,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p55_in,
            y(0) => p55_out,
            y(1 to 16 - 1) => dummy55
        );


    p56_in <= x(37) & x(39) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(72) & x(73) & x(74) & x(75) & x(76) & x(78) & x(79) & x(90) & x(91) & x(93) & x(94) & x(95) & x(102) & x(103) & x(104) & x(105) & x(106) & x(155) & x(158) & x(198) & x(199) & x(201) & x(226) & x(227) & x(249) & x(254) & x(256) & x(265) & x(268) & x(269) & x(271) & x(277) & x(280) & x(283) & x(284) & x(294) & x(295) & x(298) & x(302) & x(303) & x(305) & x(307) & x(309) & x(310) & x(311) & x(312) & x(319) & x(331) & x(332) & x(338) & x(339) & x(347) & x(361) & x(362) & x(366) & x(372) & x(376) & x(381) & x(389) & x(390) & x(401) & x(403) & x(404) & x(409) & x(418) & x(437) & x(446) & x(459) & x(464) & x(511) & x(557) & x(657) & x(664) & x(665) & x(666) & x(693) & x(694) & x(695) & x(708) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(735) & x(736) & x(748) & x(749) & x(764) & x(769) & x(770) & x(771) & x(772) & x(773) & x(774);
    y(56) <= not(p56_out);
    p56 : perceptron
        Generic map (
            WEIGHTS => "00000000000000000000000000001111111011111101111111101111101111011100011000010100101000000100000011001111111",
            SHIFT => 4,
            B => -143,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p56_in,
            y(0) => p56_out,
            y(1 to 16 - 1) => dummy56
        );


    p57_in <= x(39) & x(40) & x(44) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(73) & x(78) & x(79) & x(91) & x(93) & x(94) & x(95) & x(96) & x(104) & x(105) & x(106) & x(136) & x(157) & x(163) & x(171) & x(270) & x(277) & x(323) & x(324) & x(341) & x(342) & x(350) & x(438) & x(445) & x(472) & x(473) & x(485) & x(487) & x(500) & x(501) & x(512) & x(513) & x(514) & x(515) & x(516) & x(528) & x(529) & x(541) & x(542) & x(543) & x(556) & x(557) & x(584) & x(611) & x(612) & x(675) & x(677) & x(678) & x(679) & x(693) & x(694) & x(706) & x(708) & x(709) & x(711) & x(712) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(742) & x(743) & x(744) & x(746) & x(747) & x(748);
    y(57) <= not(p57_out);
    p57 : perceptron
        Generic map (
            WEIGHTS => "0000000000000000000000101111111111000000000000000000000011111111111111111111111",
            SHIFT => 4,
            B => -124,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p57_in,
            y(0) => p57_out,
            y(1 to 16 - 1) => dummy57
        );


    p58_in <= x(78) & x(79) & x(94) & x(104) & x(105) & x(106) & x(107) & x(153) & x(199) & x(215) & x(220) & x(221) & x(222) & x(242) & x(248) & x(249) & x(250) & x(269) & x(276) & x(277) & x(278) & x(294) & x(295) & x(322) & x(330) & x(333) & x(350) & x(361) & x(362) & x(370) & x(371) & x(373) & x(431) & x(458) & x(466) & x(473) & x(483) & x(486) & x(487) & x(488) & x(501) & x(513) & x(514) & x(515) & x(516) & x(528) & x(529) & x(530) & x(543) & x(545) & x(547) & x(554) & x(555) & x(557) & x(574) & x(584) & x(611) & x(612) & x(675) & x(676) & x(677) & x(678) & x(764) & x(765);
    y(58) <= not(p58_out);
    p58 : perceptron
        Generic map (
            WEIGHTS => "1111111100000000000000001000000011011111111111111111111111000000",
            SHIFT => 4,
            B => 25,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p58_in,
            y(0) => p58_out,
            y(1 to 16 - 1) => dummy58
        );


    p59_in <= x(104) & x(105) & x(106) & x(108) & x(192) & x(198) & x(221) & x(226) & x(248) & x(249) & x(250) & x(254) & x(263) & x(264) & x(276) & x(277) & x(282) & x(283) & x(284) & x(291) & x(292) & x(295) & x(301) & x(302) & x(303) & x(305) & x(309) & x(310) & x(311) & x(322) & x(323) & x(329) & x(330) & x(331) & x(337) & x(338) & x(339) & x(349) & x(350) & x(351) & x(357) & x(358) & x(366) & x(370) & x(377) & x(378) & x(390) & x(394) & x(398) & x(400) & x(416) & x(418) & x(446) & x(450) & x(473) & x(474) & x(485) & x(501) & x(502) & x(507) & x(513) & x(514) & x(515) & x(528) & x(529) & x(530) & x(535) & x(556) & x(557) & x(558) & x(584) & x(612) & x(647) & x(648) & x(675) & x(676) & x(677) & x(678) & x(693) & x(694) & x(695) & x(707) & x(714) & x(715) & x(716) & x(717) & x(735) & x(736) & x(737) & x(738) & x(739) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(750) & x(761) & x(764) & x(765) & x(766) & x(769) & x(770) & x(771) & x(772) & x(773) & x(774);
    y(59) <= not(p59_out);
    p59 : perceptron
        Generic map (
            WEIGHTS => "0000101011100011000001000100011000000111000111001110010000010000001000001111111110000000000000000000000000000",
            SHIFT => 4,
            B => -709,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p59_in,
            y(0) => p59_out,
            y(1 to 16 - 1) => dummy59
        );


    p60_in <= x(35) & x(36) & x(37) & x(38) & x(39) & x(40) & x(41) & x(42) & x(43) & x(44) & x(45) & x(46) & x(47) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(79) & x(80) & x(90) & x(91) & x(93) & x(94) & x(95) & x(96) & x(97) & x(98) & x(99) & x(100) & x(101) & x(102) & x(103) & x(104) & x(105) & x(106) & x(107) & x(108) & x(135) & x(150) & x(153) & x(162) & x(163) & x(164) & x(165) & x(182) & x(190) & x(191) & x(192) & x(193) & x(200) & x(219) & x(226) & x(247) & x(248) & x(249) & x(263) & x(288) & x(290) & x(291) & x(294) & x(314) & x(315) & x(316) & x(317) & x(318) & x(319) & x(386) & x(396) & x(397) & x(409) & x(418) & x(425) & x(445) & x(446) & x(450) & x(464) & x(478) & x(479) & x(492) & x(497) & x(498) & x(507) & x(515) & x(534) & x(535) & x(542) & x(543) & x(544) & x(550) & x(562) & x(563) & x(573) & x(591) & x(602) & x(619) & x(620) & x(622) & x(623) & x(647) & x(648) & x(649) & x(674) & x(675) & x(676) & x(677) & x(678) & x(679) & x(690) & x(691) & x(720) & x(721) & x(723) & x(737) & x(738) & x(739) & x(740);
    y(60) <= not(p60_out);
    p60 : perceptron
        Generic map (
            WEIGHTS => "000000000000000000000000000000000000000000000000001001111011110111111111011111101111101010010000000000000000000000000000110000000",
            SHIFT => 4,
            B => -853,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p60_in,
            y(0) => p60_out,
            y(1 to 17 - 1) => dummy60
        );


    p61_in <= x(34) & x(35) & x(36) & x(37) & x(38) & x(39) & x(40) & x(41) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(79) & x(102) & x(103) & x(104) & x(105) & x(106) & x(118) & x(148) & x(151) & x(154) & x(172) & x(173) & x(174) & x(176) & x(178) & x(180) & x(181) & x(182) & x(193) & x(199) & x(200) & x(201) & x(202) & x(214) & x(215) & x(220) & x(228) & x(248) & x(249) & x(267) & x(268) & x(269) & x(276) & x(277) & x(291) & x(292) & x(294) & x(295) & x(296) & x(297) & x(298) & x(309) & x(311) & x(317) & x(319) & x(320) & x(323) & x(324) & x(338) & x(339) & x(343) & x(344) & x(347) & x(349) & x(366) & x(386) & x(390) & x(414) & x(418) & x(422) & x(446) & x(473) & x(474) & x(487) & x(495) & x(501) & x(502) & x(507) & x(515) & x(528) & x(529) & x(530) & x(534) & x(535) & x(537) & x(542) & x(550) & x(556) & x(557) & x(558) & x(563) & x(564) & x(565) & x(566) & x(579) & x(584) & x(591) & x(593) & x(595) & x(612) & x(619) & x(620) & x(652) & x(654) & x(676) & x(677) & x(691) & x(692) & x(693) & x(694) & x(695) & x(706) & x(719) & x(720) & x(721) & x(722) & x(723) & x(769) & x(770) & x(773) & x(774);
    y(61) <= not(p61_out);
    p61 : perceptron
        Generic map (
            WEIGHTS => "0000000000000000000000000000000111111111111011111101001110000111111100011110000101011111011110111111011111111111111111111000001000001111",
            SHIFT => 4,
            B => 54,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p61_in,
            y(0) => p61_out,
            y(1 to 17 - 1) => dummy61
        );


    p62_in <= x(122) & x(171) & x(192) & x(193) & x(194) & x(220) & x(221) & x(222) & x(248) & x(249) & x(250) & x(262) & x(276) & x(277) & x(278) & x(289) & x(290) & x(291) & x(302) & x(303) & x(326) & x(329) & x(330) & x(331) & x(332) & x(356) & x(357) & x(358) & x(359) & x(397) & x(400) & x(416) & x(433) & x(434) & x(450) & x(484) & x(485) & x(486) & x(487) & x(488) & x(495) & x(506) & x(507) & x(513) & x(514) & x(515) & x(516) & x(523) & x(525) & x(534) & x(535) & x(538) & x(542) & x(550) & x(563) & x(564) & x(566) & x(591) & x(618) & x(619) & x(623) & x(647) & x(648) & x(649) & x(675) & x(676) & x(677) & x(678) & x(706) & x(707) & x(708) & x(743) & x(772);
    y(62) <= not(p62_out);
    p62 : perceptron
        Generic map (
            WEIGHTS => "1111111111101110000000000000011100100000111000011111011111111111111111100",
            SHIFT => 4,
            B => 453,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p62_in,
            y(0) => p62_out,
            y(1 to 16 - 1) => dummy62
        );


    p63_in <= x(0) & x(3) & x(4) & x(5) & x(7) & x(9) & x(11) & x(12) & x(17) & x(20) & x(22) & x(23) & x(24) & x(25) & x(27) & x(28) & x(30) & x(31) & x(32) & x(35) & x(44) & x(53) & x(54) & x(55) & x(56) & x(58) & x(59) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(79) & x(80) & x(82) & x(83) & x(85) & x(88) & x(93) & x(94) & x(95) & x(96) & x(97) & x(101) & x(102) & x(103) & x(104) & x(105) & x(106) & x(107) & x(108) & x(110) & x(111) & x(112) & x(113) & x(118) & x(133) & x(135) & x(139) & x(148) & x(155) & x(165) & x(169) & x(171) & x(172) & x(173) & x(176) & x(190) & x(192) & x(196) & x(197) & x(199) & x(200) & x(201) & x(221) & x(227) & x(228) & x(248) & x(249) & x(256) & x(277) & x(283) & x(284) & x(304) & x(309) & x(310) & x(311) & x(312) & x(330) & x(332) & x(333) & x(337) & x(338) & x(339) & x(342) & x(346) & x(350) & x(361) & x(362) & x(366) & x(367) & x(369) & x(370) & x(371) & x(372) & x(374) & x(387) & x(389) & x(390) & x(392) & x(396) & x(397) & x(398) & x(399) & x(400) & x(401) & x(410) & x(417) & x(422) & x(428) & x(430) & x(431) & x(434) & x(445) & x(448) & x(450) & x(451) & x(473) & x(474) & x(478) & x(479) & x(502) & x(504) & x(507) & x(515) & x(532) & x(534) & x(535) & x(557) & x(560) & x(562) & x(563) & x(587) & x(588) & x(591) & x(615) & x(616) & x(618) & x(619) & x(620) & x(644) & x(647) & x(665) & x(671) & x(673) & x(692) & x(693) & x(694) & x(698) & x(700) & x(702) & x(719) & x(721) & x(722) & x(725) & x(726) & x(727) & x(730) & x(731) & x(748) & x(753) & x(754) & x(757) & x(758) & x(764) & x(765) & x(766) & x(768) & x(769) & x(770) & x(771) & x(772) & x(773) & x(774) & x(780) & x(781);
    y(63) <= not(p63_out);
    p63 : perceptron
        Generic map (
            WEIGHTS => "0000000000000000000110000001111111111111100001111111111111000010001100111100011110110010111111111111100111110000001100000001110001101111111011011101100100111010000000000000000000000111111111100",
            SHIFT => 4,
            B => 64,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p63_in,
            y(0) => p63_out,
            y(1 to 17 - 1) => dummy63
        );


    p64_in <= x(36) & x(37) & x(38) & x(39) & x(40) & x(41) & x(44) & x(45) & x(46) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(79) & x(90) & x(91) & x(92) & x(93) & x(94) & x(103) & x(104) & x(105) & x(106) & x(126) & x(127) & x(135) & x(164) & x(165) & x(166) & x(191) & x(192) & x(193) & x(194) & x(198) & x(207) & x(208) & x(209) & x(219) & x(220) & x(221) & x(222) & x(234) & x(235) & x(245) & x(247) & x(248) & x(249) & x(250) & x(254) & x(276) & x(277) & x(278) & x(288) & x(295) & x(297) & x(298) & x(299) & x(300) & x(302) & x(303) & x(304) & x(305) & x(306) & x(315) & x(320) & x(327) & x(328) & x(329) & x(330) & x(331) & x(332) & x(339) & x(340) & x(342) & x(343) & x(347) & x(348) & x(357) & x(358) & x(359) & x(360) & x(376) & x(377) & x(380) & x(381) & x(388) & x(404) & x(408) & x(425) & x(446) & x(453) & x(454) & x(456) & x(474) & x(479) & x(481) & x(483) & x(502) & x(507) & x(517) & x(518) & x(529) & x(544) & x(545) & x(546) & x(557) & x(584) & x(611) & x(612) & x(626) & x(633) & x(652) & x(653) & x(654) & x(655) & x(656) & x(657) & x(660) & x(677) & x(679) & x(681) & x(682) & x(684) & x(685) & x(706) & x(707) & x(708) & x(709) & x(710) & x(711) & x(712) & x(715) & x(720) & x(737) & x(739) & x(742) & x(743) & x(744) & x(746) & x(761) & x(764) & x(765) & x(766) & x(770) & x(773) & x(774);
    y(64) <= not(p64_out);
    p64 : perceptron
        Generic map (
            WEIGHTS => "000000000000000000000000000000000000110000000000000000000000000000111111110000111111000000111100000001111110111011111111110000000000000000000000000000000000000",
            SHIFT => 3,
            B => -812,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p64_in,
            y(0) => p64_out,
            y(1 to 16 - 1) => dummy64
        );


    p65_in <= x(35) & x(41) & x(63) & x(64) & x(68) & x(79) & x(105) & x(108) & x(135) & x(163) & x(164) & x(191) & x(192) & x(193) & x(194) & x(195) & x(220) & x(221) & x(222) & x(248) & x(249) & x(250) & x(276) & x(277) & x(278) & x(303) & x(305) & x(306) & x(310) & x(329) & x(330) & x(331) & x(332) & x(333) & x(334) & x(338) & x(339) & x(346) & x(347) & x(349) & x(358) & x(359) & x(360) & x(366) & x(374) & x(375) & x(376) & x(377) & x(378) & x(388) & x(450) & x(479) & x(507) & x(514) & x(515) & x(535) & x(542) & x(543) & x(544) & x(591) & x(648) & x(655) & x(656) & x(657) & x(675) & x(677);
    y(65) <= not(p65_out);
    p65 : perceptron
        Generic map (
            WEIGHTS => "111111110000000000000000010011111001100011110000010001101110000000",
            SHIFT => 4,
            B => -169,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p65_in,
            y(0) => p65_out,
            y(1 to 16 - 1) => dummy65
        );


    p66_in <= x(34) & x(35) & x(36) & x(37) & x(38) & x(39) & x(40) & x(41) & x(42) & x(43) & x(44) & x(45) & x(46) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(79) & x(80) & x(90) & x(91) & x(92) & x(93) & x(94) & x(95) & x(96) & x(97) & x(98) & x(99) & x(100) & x(101) & x(102) & x(103) & x(104) & x(105) & x(106) & x(107) & x(108) & x(135) & x(136) & x(163) & x(164) & x(191) & x(192) & x(303) & x(304) & x(321) & x(323) & x(324) & x(329) & x(330) & x(331) & x(332) & x(348) & x(349) & x(358) & x(359) & x(368) & x(369) & x(370) & x(376) & x(387) & x(388) & x(396) & x(397) & x(398) & x(418) & x(425) & x(426) & x(446) & x(451) & x(453) & x(475) & x(479) & x(487) & x(488) & x(501) & x(507) & x(513) & x(514) & x(515) & x(516) & x(528) & x(529) & x(530) & x(534) & x(541) & x(542) & x(543) & x(544) & x(556) & x(557) & x(570) & x(571) & x(584) & x(591) & x(647);
    y(66) <= not(p66_out);
    p66 : perceptron
        Generic map (
            WEIGHTS => "11111111111111111111111111111111111111111111111111100000011100111111110001110000000100111011111000111110011011",
            SHIFT => 4,
            B => 686,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p66_in,
            y(0) => p66_out,
            y(1 to 16 - 1) => dummy66
        );


    p67_in <= x(63) & x(166) & x(171) & x(192) & x(193) & x(198) & x(199) & x(219) & x(220) & x(239) & x(247) & x(248) & x(249) & x(266) & x(267) & x(276) & x(277) & x(294) & x(295) & x(296) & x(309) & x(319) & x(322) & x(323) & x(339) & x(347) & x(348) & x(361) & x(362) & x(366) & x(375) & x(376) & x(379) & x(390) & x(418) & x(422) & x(474) & x(485) & x(486) & x(513) & x(514) & x(542) & x(543) & x(665) & x(676) & x(677) & x(693) & x(694) & x(764) & x(773) & x(774);
    y(67) <= not(p67_out);
    p67 : perceptron
        Generic map (
            WEIGHTS => "001001100100011001111011100111001111111111101100111",
            SHIFT => 4,
            B => 157,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p67_in,
            y(0) => p67_out,
            y(1 to 15 - 1) => dummy67
        );


    p68_in <= x(64) & x(65) & x(67) & x(68) & x(70) & x(72) & x(73) & x(74) & x(75) & x(76) & x(78) & x(79) & x(104) & x(105) & x(106) & x(151) & x(152) & x(179) & x(180) & x(182) & x(186) & x(199) & x(211) & x(213) & x(239) & x(248) & x(249) & x(250) & x(271) & x(272) & x(275) & x(276) & x(299) & x(303) & x(304) & x(307) & x(332) & x(361) & x(362) & x(366) & x(390) & x(401) & x(423) & x(434) & x(462) & x(489) & x(517) & x(518) & x(574) & x(622) & x(657) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(748) & x(749) & x(750);
    y(68) <= not(p68_out);
    p68 : perceptron
        Generic map (
            WEIGHTS => "00000000000000011111111111111111111111111000000001111111111111111111",
            SHIFT => 4,
            B => 364,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p68_in,
            y(0) => p68_out,
            y(1 to 16 - 1) => dummy68
        );


    p69_in <= x(64) & x(67) & x(68) & x(70) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(79) & x(102) & x(103) & x(104) & x(105) & x(106) & x(107) & x(126) & x(127) & x(133) & x(163) & x(188) & x(189) & x(190) & x(201) & x(221) & x(235) & x(243) & x(248) & x(249) & x(250) & x(267) & x(269) & x(276) & x(277) & x(278) & x(283) & x(284) & x(307) & x(312) & x(333) & x(338) & x(339) & x(357) & x(358) & x(359) & x(361) & x(362) & x(366) & x(367) & x(389) & x(390) & x(406) & x(418) & x(432) & x(433) & x(434) & x(458) & x(467) & x(486) & x(487) & x(488) & x(490) & x(514) & x(515) & x(516) & x(518) & x(666) & x(675) & x(677) & x(721) & x(748) & x(769) & x(770) & x(773);
    y(69) <= not(p69_out);
    p69 : perceptron
        Generic map (
            WEIGHTS => "0000000000000000000011111111111111111111111100011111101000010000000001100111",
            SHIFT => 4,
            B => 52,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p69_in,
            y(0) => p69_out,
            y(1 to 16 - 1) => dummy69
        );


    p70_in <= x(35) & x(43) & x(75) & x(97) & x(108) & x(164) & x(165) & x(166) & x(182) & x(183) & x(191) & x(192) & x(193) & x(209) & x(210) & x(211) & x(212) & x(219) & x(220) & x(221) & x(237) & x(238) & x(239) & x(240) & x(247) & x(248) & x(249) & x(266) & x(267) & x(268) & x(276) & x(277) & x(294) & x(295) & x(305) & x(306) & x(320) & x(329) & x(333) & x(334) & x(338) & x(347) & x(348) & x(349) & x(366) & x(376) & x(377) & x(433) & x(450) & x(460) & x(474) & x(501) & x(507) & x(514) & x(515) & x(529) & x(534) & x(535) & x(557) & x(563) & x(591) & x(618) & x(638) & x(647) & x(648) & x(675) & x(703) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(732) & x(738) & x(739) & x(740) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(748) & x(749);
    y(70) <= not(p70_out);
    p70 : perceptron
        Generic map (
            WEIGHTS => "10011000110001111000111100011100110001001000100000110111001000100001111111111111111111",
            SHIFT => 4,
            B => -45,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p70_in,
            y(0) => p70_out,
            y(1 to 16 - 1) => dummy70
        );


    p71_in <= x(35) & x(37) & x(38) & x(40) & x(41) & x(62) & x(63) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(210) & x(218) & x(219) & x(238) & x(266) & x(267) & x(275) & x(277) & x(294) & x(295) & x(302) & x(303) & x(322) & x(323) & x(330) & x(331) & x(342) & x(405) & x(424) & x(425) & x(432) & x(433) & x(434) & x(446) & x(453) & x(460) & x(461) & x(473) & x(474) & x(484) & x(485) & x(487) & x(488) & x(500) & x(501) & x(502) & x(512) & x(513) & x(514) & x(515) & x(516) & x(528) & x(529) & x(556) & x(557) & x(558) & x(584) & x(648) & x(675) & x(676) & x(677) & x(678) & x(694) & x(695) & x(706) & x(708) & x(709) & x(710) & x(711) & x(712) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(737) & x(739) & x(740) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(748) & x(749) & x(764) & x(765) & x(766);
    y(71) <= not(p71_out);
    p71 : perceptron
        Generic map (
            WEIGHTS => "000000000000001100010001100110111111111111111111111111111111000000000000000000000000000000000000",
            SHIFT => 4,
            B => -358,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p71_in,
            y(0) => p71_out,
            y(1 to 16 - 1) => dummy71
        );


    p72_in <= x(67) & x(68) & x(69) & x(97) & x(99) & x(108) & x(157) & x(191) & x(192) & x(193) & x(210) & x(212) & x(219) & x(220) & x(237) & x(248) & x(266) & x(294) & x(334) & x(348) & x(349) & x(366) & x(374) & x(377) & x(432) & x(433) & x(473) & x(515) & x(529) & x(535) & x(543) & x(557) & x(563) & x(584) & x(591) & x(605) & x(619) & x(647) & x(667) & x(708) & x(709) & x(711) & x(712) & x(713) & x(715) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(736) & x(737) & x(738) & x(739) & x(740) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(748) & x(749) & x(764);
    y(72) <= not(p72_out);
    p72 : perceptron
        Generic map (
            WEIGHTS => "00000011110011010011101111101101111111100000000000000000000000000000",
            SHIFT => 5,
            B => -394,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p72_in,
            y(0) => p72_out,
            y(1 to 17 - 1) => dummy72
        );


    p73_in <= x(132) & x(133) & x(166) & x(193) & x(220) & x(221) & x(247) & x(248) & x(249) & x(250) & x(269) & x(275) & x(276) & x(277) & x(278) & x(303) & x(304) & x(305) & x(306) & x(307) & x(320) & x(321) & x(333) & x(334) & x(348) & x(349) & x(361) & x(362) & x(367) & x(376) & x(380) & x(389) & x(390) & x(407) & x(408) & x(414) & x(432) & x(433) & x(450) & x(479) & x(487) & x(514) & x(535) & x(656) & x(666);
    y(73) <= not(p73_out);
    p73 : perceptron
        Generic map (
            WEIGHTS => "110000000010000000000000000000000000000000001",
            SHIFT => 5,
            B => -731,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p73_in,
            y(0) => p73_out,
            y(1 to 16 - 1) => dummy73
        );


    p74_in <= x(34) & x(35) & x(37) & x(39) & x(40) & x(41) & x(62) & x(63) & x(64) & x(66) & x(68) & x(69) & x(75) & x(109) & x(118) & x(146) & x(147) & x(172) & x(173) & x(174) & x(248) & x(266) & x(276) & x(295) & x(296) & x(297) & x(305) & x(320) & x(323) & x(348) & x(410) & x(414) & x(416) & x(418) & x(437) & x(444) & x(446) & x(450) & x(457) & x(459) & x(473) & x(474) & x(475) & x(479) & x(486) & x(487) & x(501) & x(502) & x(507) & x(513) & x(514) & x(529) & x(530) & x(534) & x(535) & x(542) & x(543) & x(544) & x(557) & x(558) & x(562) & x(563) & x(572) & x(584) & x(585) & x(591) & x(592) & x(612) & x(618) & x(619) & x(620) & x(647) & x(648) & x(676) & x(677) & x(709) & x(710) & x(711);
    y(74) <= not(p74_out);
    p74 : perceptron
        Generic map (
            WEIGHTS => "111111111111100000001010000101011001001100001100011000011100001000000000000000",
            SHIFT => 4,
            B => -370,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p74_in,
            y(0) => p74_out,
            y(1 to 16 - 1) => dummy74
        );


    p75_in <= x(37) & x(40) & x(41) & x(63) & x(64) & x(68) & x(72) & x(73) & x(74) & x(75) & x(78) & x(79) & x(103) & x(104) & x(105) & x(106) & x(107) & x(133) & x(189) & x(190) & x(198) & x(226) & x(248) & x(249) & x(250) & x(254) & x(266) & x(276) & x(277) & x(309) & x(310) & x(338) & x(339) & x(352) & x(362) & x(366) & x(377) & x(378) & x(381) & x(390) & x(394) & x(405) & x(409) & x(418) & x(431) & x(434) & x(436) & x(446) & x(450) & x(474) & x(478) & x(501) & x(502) & x(506) & x(507) & x(534) & x(535) & x(544) & x(563) & x(583) & x(591) & x(619) & x(620) & x(647) & x(648) & x(649) & x(675) & x(676) & x(693) & x(736) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(750) & x(764) & x(765) & x(766) & x(769) & x(770) & x(772) & x(773) & x(774);
    y(75) <= not(p75_out);
    p75 : perceptron
        Generic map (
            WEIGHTS => "00000000000000000111111111111111101100011001000101011000010100000000011111111111111111",
            SHIFT => 5,
            B => 227,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p75_in,
            y(0) => p75_out,
            y(1 to 17 - 1) => dummy75
        );


    p76_in <= x(76) & x(96) & x(101) & x(102) & x(103) & x(106) & x(108) & x(133) & x(163) & x(164) & x(165) & x(191) & x(192) & x(200) & x(219) & x(220) & x(221) & x(247) & x(248) & x(249) & x(275) & x(277) & x(301) & x(302) & x(303) & x(304) & x(305) & x(320) & x(323) & x(327) & x(329) & x(330) & x(331) & x(332) & x(333) & x(338) & x(344) & x(347) & x(358) & x(361) & x(362) & x(371) & x(390) & x(418) & x(445) & x(446) & x(473) & x(474) & x(475) & x(479) & x(502) & x(507) & x(529) & x(535) & x(557) & x(563) & x(591) & x(619) & x(647) & x(715) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(723) & x(740) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(748) & x(769) & x(770);
    y(76) <= not(p76_out);
    p76 : perceptron
        Generic map (
            WEIGHTS => "000000011111101111111100000100000000110001000000000000000000000000000000000000",
            SHIFT => 5,
            B => -1343,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p76_in,
            y(0) => p76_out,
            y(1 to 17 - 1) => dummy76
        );


    p77_in <= x(40) & x(41) & x(73) & x(74) & x(198) & x(226) & x(254) & x(282) & x(309) & x(310) & x(311) & x(338) & x(339) & x(340) & x(349) & x(359) & x(360) & x(366) & x(367) & x(368) & x(387) & x(388) & x(394) & x(397) & x(400) & x(413) & x(414) & x(415) & x(416) & x(418) & x(425) & x(443) & x(444) & x(446) & x(450) & x(473) & x(474) & x(501) & x(502) & x(506) & x(528) & x(529) & x(530) & x(556) & x(557) & x(558) & x(583) & x(584) & x(611) & x(612) & x(640) & x(647) & x(675) & x(707) & x(708) & x(709) & x(710) & x(711) & x(712) & x(713) & x(714) & x(715) & x(716) & x(717) & x(718) & x(719) & x(735) & x(736) & x(737) & x(738) & x(739) & x(740) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(748) & x(750) & x(764) & x(765) & x(766) & x(769) & x(770) & x(771) & x(772) & x(773) & x(774) & x(775);
    y(77) <= not(p77_out);
    p77 : perceptron
        Generic map (
            WEIGHTS => "0000111111111100011100100000010001011110111111111110011111111111111111111111111111111111111",
            SHIFT => 5,
            B => 1297,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p77_in,
            y(0) => p77_out,
            y(1 to 17 - 1) => dummy77
        );


    p78_in <= x(67) & x(68) & x(69) & x(152) & x(179) & x(180) & x(182) & x(183) & x(185) & x(193) & x(220) & x(221) & x(248) & x(249) & x(250) & x(276) & x(293) & x(297) & x(304) & x(306) & x(307) & x(320) & x(325) & x(331) & x(332) & x(334) & x(348) & x(349) & x(354) & x(360) & x(361) & x(362) & x(376) & x(381) & x(388) & x(389) & x(390) & x(411) & x(437) & x(444) & x(450) & x(464) & x(469) & x(491) & x(506) & x(517) & x(523) & x(529) & x(530) & x(534) & x(542) & x(557) & x(566) & x(568) & x(569) & x(578) & x(584) & x(597) & x(622) & x(647) & x(653) & x(655) & x(656) & x(657) & x(658) & x(666) & x(674) & x(675) & x(712) & x(737) & x(739) & x(742) & x(761);
    y(78) <= not(p78_out);
    p78 : perceptron
        Generic map (
            WEIGHTS => "0000000000000000110000100000100001000110010101011001000010000000010011111",
            SHIFT => 4,
            B => -372,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p78_in,
            y(0) => p78_out,
            y(1 to 16 - 1) => dummy78
        );


    p79_in <= x(78) & x(105) & x(106) & x(107) & x(108) & x(162) & x(166) & x(192) & x(194) & x(195) & x(219) & x(220) & x(221) & x(222) & x(247) & x(248) & x(249) & x(250) & x(276) & x(277) & x(278) & x(289) & x(297) & x(298) & x(299) & x(305) & x(306) & x(323) & x(324) & x(325) & x(326) & x(327) & x(328) & x(329) & x(330) & x(331) & x(350) & x(351) & x(353) & x(358) & x(362) & x(377) & x(378) & x(381) & x(390) & x(408) & x(409) & x(416) & x(418) & x(433) & x(436) & x(437) & x(464) & x(474) & x(514) & x(515) & x(638) & x(681) & x(682) & x(690) & x(692) & x(693) & x(719) & x(720) & x(721) & x(722) & x(748) & x(764) & x(765);
    y(79) <= not(p79_out);
    p79 : perceptron
        Generic map (
            WEIGHTS => "111110000000000000000011100111111111111101110110011110110111111111100",
            SHIFT => 4,
            B => -26,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p79_in,
            y(0) => p79_out,
            y(1 to 16 - 1) => dummy79
        );


    p80_in <= x(96) & x(104) & x(105) & x(106) & x(156) & x(157) & x(210) & x(211) & x(238) & x(248) & x(249) & x(250) & x(266) & x(267) & x(276) & x(277) & x(294) & x(295) & x(305) & x(311) & x(322) & x(323) & x(333) & x(349) & x(350) & x(351) & x(360) & x(377) & x(378) & x(432) & x(473) & x(485) & x(501) & x(502) & x(512) & x(528) & x(529) & x(530) & x(556) & x(557) & x(558) & x(584) & x(611) & x(612) & x(638) & x(692) & x(693) & x(694) & x(695) & x(709) & x(712) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(724) & x(742) & x(745) & x(746) & x(747) & x(748) & x(749);
    y(80) <= not(p80_out);
    p80 : perceptron
        Generic map (
            WEIGHTS => "111111000000000000010000001001111111111111111000000000000000000000",
            SHIFT => 4,
            B => -180,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p80_in,
            y(0) => p80_out,
            y(1 to 16 - 1) => dummy80
        );


    p81_in <= x(91) & x(93) & x(94) & x(95) & x(96) & x(100) & x(102) & x(125) & x(147) & x(148) & x(150) & x(151) & x(176) & x(178) & x(179) & x(198) & x(260) & x(287) & x(289) & x(291) & x(316) & x(317) & x(322) & x(327) & x(333) & x(342) & x(343) & x(344) & x(350) & x(354) & x(355) & x(361) & x(376) & x(378) & x(400) & x(401) & x(403) & x(406) & x(428) & x(431) & x(434) & x(450) & x(472) & x(473) & x(474) & x(501) & x(502) & x(508) & x(521) & x(522) & x(526) & x(528) & x(529) & x(535) & x(536) & x(549) & x(556) & x(557) & x(558) & x(563) & x(564) & x(565) & x(578) & x(579) & x(580) & x(584) & x(585) & x(586) & x(591) & x(592) & x(611) & x(612) & x(619) & x(620) & x(622) & x(638) & x(647) & x(649) & x(650) & x(657) & x(675) & x(676) & x(677) & x(690) & x(691) & x(692) & x(693) & x(694) & x(695) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(742) & x(746) & x(747) & x(748);
    y(81) <= not(p81_out);
    p81 : perceptron
        Generic map (
            WEIGHTS => "111111111111111000000000000000001011101101111111111111111111111111111111111111101110000000000000000",
            SHIFT => 4,
            B => 366,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p81_in,
            y(0) => p81_out,
            y(1 to 16 - 1) => dummy81
        );


    p82_in <= x(3) & x(21) & x(22) & x(25) & x(26) & x(30) & x(35) & x(57) & x(63) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(79) & x(82) & x(96) & x(106) & x(108) & x(113) & x(118) & x(153) & x(154) & x(168) & x(171) & x(172) & x(173) & x(200) & x(248) & x(303) & x(304) & x(305) & x(322) & x(333) & x(338) & x(339) & x(350) & x(361) & x(362) & x(366) & x(367) & x(370) & x(371) & x(377) & x(389) & x(390) & x(396) & x(397) & x(398) & x(399) & x(401) & x(405) & x(406) & x(413) & x(427) & x(428) & x(429) & x(430) & x(433) & x(434) & x(445) & x(450) & x(451) & x(473) & x(474) & x(478) & x(479) & x(507) & x(534) & x(535) & x(562) & x(563) & x(574) & x(591) & x(607) & x(615) & x(618) & x(619) & x(624) & x(643) & x(647) & x(648) & x(653) & x(654) & x(656) & x(658) & x(725) & x(727) & x(729) & x(730) & x(754) & x(756) & x(770) & x(771) & x(773) & x(774) & x(780);
    y(82) <= not(p82_out);
    p82 : perceptron
        Generic map (
            WEIGHTS => "00000010111111110111011101111111111111111100111000001100000111111111111110110111011111100000011110",
            SHIFT => 4,
            B => 38,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p82_in,
            y(0) => p82_out,
            y(1 to 16 - 1) => dummy82
        );


    p83_in <= x(63) & x(64) & x(79) & x(91) & x(136) & x(164) & x(165) & x(166) & x(171) & x(172) & x(191) & x(192) & x(193) & x(194) & x(197) & x(220) & x(221) & x(222) & x(248) & x(249) & x(250) & x(266) & x(276) & x(277) & x(278) & x(296) & x(297) & x(305) & x(306) & x(307) & x(322) & x(323) & x(328) & x(329) & x(333) & x(334) & x(338) & x(346) & x(348) & x(349) & x(350) & x(351) & x(358) & x(359) & x(361) & x(362) & x(377) & x(378) & x(406) & x(423) & x(433) & x(434) & x(450) & x(454) & x(461) & x(473) & x(474) & x(478) & x(479) & x(501) & x(502) & x(506) & x(507) & x(511) & x(512) & x(514) & x(528) & x(529) & x(530) & x(534) & x(535) & x(543) & x(546) & x(556) & x(557) & x(558) & x(563) & x(584) & x(591) & x(600) & x(611) & x(612) & x(618) & x(638) & x(639) & x(646) & x(647) & x(648) & x(649) & x(658) & x(674) & x(675) & x(676) & x(677) & x(678) & x(679) & x(716) & x(720) & x(732) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747);
    y(83) <= not(p83_out);
    p83 : perceptron
        Generic map (
            WEIGHTS => "0000111111111111111110111001111100110111110011111111101001100110000001100000101000100111111111110100000000",
            SHIFT => 4,
            B => 238,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p83_in,
            y(0) => p83_out,
            y(1 to 16 - 1) => dummy83
        );


    p84_in <= x(37) & x(40) & x(41) & x(45) & x(46) & x(48) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(103) & x(104) & x(105) & x(106) & x(135) & x(136) & x(163) & x(164) & x(165) & x(166) & x(191) & x(192) & x(193) & x(194) & x(199) & x(219) & x(220) & x(221) & x(222) & x(227) & x(247) & x(248) & x(249) & x(250) & x(254) & x(276) & x(277) & x(278) & x(298) & x(299) & x(300) & x(301) & x(302) & x(303) & x(304) & x(305) & x(306) & x(320) & x(326) & x(327) & x(328) & x(329) & x(330) & x(331) & x(332) & x(347) & x(348) & x(357) & x(358) & x(359) & x(360) & x(390) & x(418) & x(425) & x(446) & x(450) & x(453) & x(454) & x(473) & x(474) & x(481) & x(485) & x(487) & x(501) & x(502) & x(512) & x(513) & x(514) & x(515) & x(529) & x(542) & x(543) & x(556) & x(557) & x(584) & x(612) & x(639) & x(640) & x(648) & x(675) & x(676) & x(677) & x(678) & x(679) & x(706) & x(707) & x(708) & x(709) & x(711) & x(712) & x(718) & x(720) & x(734) & x(735) & x(736) & x(737) & x(739) & x(742) & x(743) & x(761) & x(764) & x(765) & x(766) & x(769) & x(770) & x(771) & x(773);
    y(84) <= not(p84_out);
    p84 : perceptron
        Generic map (
            WEIGHTS => "0000000000000000000000000000000000000000000000000001111111000111111100111111110111111111111111111111100000000000011000000000000000",
            SHIFT => 4,
            B => -708,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p84_in,
            y(0) => p84_out,
            y(1 to 17 - 1) => dummy84
        );


    p85_in <= x(75) & x(99) & x(100) & x(101) & x(102) & x(103) & x(135) & x(163) & x(171) & x(172) & x(182) & x(183) & x(184) & x(192) & x(195) & x(197) & x(199) & x(200) & x(210) & x(211) & x(212) & x(220) & x(221) & x(222) & x(227) & x(228) & x(238) & x(239) & x(249) & x(255) & x(256) & x(277) & x(283) & x(294) & x(295) & x(302) & x(303) & x(305) & x(310) & x(311) & x(312) & x(322) & x(323) & x(324) & x(329) & x(330) & x(331) & x(333) & x(357) & x(358) & x(359) & x(360) & x(366) & x(422) & x(423) & x(450) & x(478) & x(479) & x(507) & x(513) & x(514) & x(515) & x(534) & x(535) & x(542) & x(563) & x(648) & x(675) & x(676) & x(677) & x(678) & x(679) & x(705) & x(706) & x(707) & x(708) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(735) & x(736) & x(747) & x(748) & x(749) & x(764) & x(769) & x(770) & x(773) & x(774);
    y(85) <= not(p85_out);
    p85 : perceptron
        Generic map (
            WEIGHTS => "000000000011100000111000001100000001100000001110111100000001110010000000000011111110011100000",
            SHIFT => 4,
            B => -687,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p85_in,
            y(0) => p85_out,
            y(1 to 16 - 1) => dummy85
        );


    p86_in <= x(64) & x(65) & x(66) & x(108) & x(133) & x(135) & x(146) & x(147) & x(162) & x(165) & x(166) & x(171) & x(172) & x(173) & x(174) & x(191) & x(192) & x(193) & x(197) & x(199) & x(200) & x(201) & x(202) & x(219) & x(220) & x(221) & x(222) & x(228) & x(247) & x(248) & x(249) & x(250) & x(261) & x(267) & x(276) & x(277) & x(290) & x(291) & x(295) & x(296) & x(297) & x(298) & x(299) & x(302) & x(304) & x(309) & x(320) & x(323) & x(326) & x(327) & x(330) & x(331) & x(332) & x(334) & x(360) & x(361) & x(366) & x(390) & x(450) & x(474) & x(478) & x(479) & x(489) & x(490) & x(502) & x(506) & x(507) & x(516) & x(534) & x(535) & x(557) & x(562) & x(563) & x(564) & x(591) & x(618) & x(619) & x(646) & x(647) & x(648) & x(675) & x(676) & x(677) & x(747) & x(750);
    y(86) <= not(p86_out);
    p86 : perceptron
        Generic map (
            WEIGHTS => "1110110011100001110000011110111110111100000000100000010000000011000100000000000000000",
            SHIFT => 5,
            B => -604,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p86_in,
            y(0) => p86_out,
            y(1 to 17 - 1) => dummy86
        );


    p87_in <= x(37) & x(38) & x(39) & x(40) & x(41) & x(43) & x(45) & x(46) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(79) & x(102) & x(103) & x(104) & x(105) & x(106) & x(108) & x(133) & x(164) & x(183) & x(191) & x(192) & x(193) & x(210) & x(211) & x(219) & x(220) & x(221) & x(238) & x(239) & x(240) & x(248) & x(249) & x(268) & x(276) & x(277) & x(296) & x(297) & x(298) & x(301) & x(302) & x(303) & x(305) & x(320) & x(327) & x(328) & x(329) & x(330) & x(331) & x(332) & x(338) & x(348) & x(349) & x(360) & x(390) & x(414) & x(418) & x(446) & x(473) & x(474) & x(501) & x(502) & x(528) & x(529) & x(556) & x(557) & x(558) & x(584) & x(612) & x(619) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(732) & x(736) & x(737) & x(738) & x(739) & x(740) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(748) & x(749);
    y(87) <= not(p87_out);
    p87 : perceptron
        Generic map (
            WEIGHTS => "1111111111111111111111111111111011011100111000110110000001100000001100100000000000000000000000000000000000",
            SHIFT => 4,
            B => -11,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p87_in,
            y(0) => p87_out,
            y(1 to 16 - 1) => dummy87
        );


    p88_in <= x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(91) & x(92) & x(93) & x(104) & x(105) & x(106) & x(107) & x(145) & x(194) & x(221) & x(222) & x(228) & x(248) & x(249) & x(250) & x(277) & x(278) & x(299) & x(301) & x(302) & x(303) & x(305) & x(320) & x(326) & x(327) & x(328) & x(329) & x(330) & x(331) & x(332) & x(356) & x(357) & x(358) & x(359) & x(360) & x(385) & x(386) & x(387) & x(388) & x(390) & x(414) & x(415) & x(418) & x(446) & x(473) & x(474) & x(484) & x(485) & x(500) & x(501) & x(502) & x(513) & x(514) & x(515) & x(528) & x(529) & x(556) & x(557) & x(584) & x(611) & x(612) & x(638) & x(640) & x(666) & x(690);
    y(88) <= not(p88_out);
    p88 : perceptron
        Generic map (
            WEIGHTS => "000000011100000111011111000010000000000000000010011110011100011111111110",
            SHIFT => 4,
            B => -50,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p88_in,
            y(0) => p88_out,
            y(1 to 16 - 1) => dummy88
        );


    p89_in <= x(37) & x(39) & x(41) & x(63) & x(64) & x(65) & x(66) & x(68) & x(69) & x(70) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(79) & x(103) & x(104) & x(105) & x(106) & x(107) & x(157) & x(198) & x(226) & x(227) & x(250) & x(254) & x(255) & x(256) & x(267) & x(268) & x(269) & x(282) & x(283) & x(284) & x(285) & x(294) & x(295) & x(309) & x(310) & x(311) & x(312) & x(318) & x(338) & x(339) & x(346) & x(349) & x(353) & x(358) & x(359) & x(362) & x(366) & x(367) & x(373) & x(374) & x(376) & x(377) & x(378) & x(381) & x(382) & x(386) & x(387) & x(390) & x(404) & x(409) & x(418) & x(431) & x(432) & x(433) & x(436) & x(437) & x(446) & x(460) & x(464) & x(473) & x(474) & x(478) & x(486) & x(487) & x(488) & x(500) & x(501) & x(502) & x(506) & x(509) & x(515) & x(528) & x(529) & x(556) & x(557) & x(569) & x(570) & x(571) & x(584) & x(597) & x(638) & x(690) & x(691) & x(692) & x(693) & x(694) & x(695) & x(696) & x(704) & x(706) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(735) & x(736) & x(737) & x(743) & x(744) & x(748) & x(749) & x(764) & x(765) & x(766) & x(769) & x(770) & x(771) & x(772) & x(773) & x(774);
    y(89) <= not(p89_out);
    p89 : perceptron
        Generic map (
            WEIGHTS => "111111111111111111111110000000000000000000001001111100011111111101101111101100111100010100000000001111111001111110000011000000000",
            SHIFT => 4,
            B => -70,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p89_in,
            y(0) => p89_out,
            y(1 to 17 - 1) => dummy89
        );


    p90_in <= x(35) & x(37) & x(38) & x(39) & x(40) & x(41) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(79) & x(90) & x(91) & x(92) & x(93) & x(94) & x(95) & x(96) & x(97) & x(98) & x(99) & x(100) & x(101) & x(102) & x(103) & x(104) & x(105) & x(106) & x(107) & x(108) & x(163) & x(241) & x(242) & x(243) & x(248) & x(268) & x(295) & x(330) & x(338) & x(369) & x(396) & x(397) & x(398) & x(400) & x(425) & x(433) & x(434) & x(445) & x(454) & x(455) & x(462) & x(473) & x(487) & x(513) & x(514) & x(515) & x(516) & x(519) & x(541) & x(542) & x(543) & x(544) & x(584) & x(636) & x(640) & x(679) & x(680) & x(709) & x(710) & x(737) & x(738) & x(743);
    y(90) <= not(p90_out);
    p90 : perceptron
        Generic map (
            WEIGHTS => "000000000000000000000000000000000000000000111111100111111000000000000000000001111000",
            SHIFT => 4,
            B => -597,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p90_in,
            y(0) => p90_out,
            y(1 to 16 - 1) => dummy90
        );


    p91_in <= x(35) & x(37) & x(39) & x(40) & x(41) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(77) & x(78) & x(92) & x(104) & x(105) & x(106) & x(109) & x(125) & x(147) & x(148) & x(152) & x(153) & x(154) & x(155) & x(162) & x(165) & x(166) & x(171) & x(172) & x(176) & x(182) & x(190) & x(191) & x(192) & x(193) & x(198) & x(200) & x(210) & x(219) & x(221) & x(226) & x(248) & x(249) & x(254) & x(260) & x(267) & x(276) & x(277) & x(289) & x(292) & x(294) & x(295) & x(296) & x(297) & x(299) & x(300) & x(301) & x(302) & x(303) & x(317) & x(320) & x(323) & x(327) & x(332) & x(342) & x(343) & x(344) & x(347) & x(348) & x(370) & x(371) & x(373) & x(374) & x(378) & x(401) & x(402) & x(418) & x(446) & x(450) & x(473) & x(474) & x(475) & x(479) & x(501) & x(502) & x(507) & x(529) & x(534) & x(535) & x(557) & x(562) & x(563) & x(564) & x(566) & x(584) & x(591) & x(594) & x(601) & x(612) & x(618) & x(619) & x(620) & x(623) & x(647) & x(648) & x(677) & x(721) & x(723) & x(748);
    y(91) <= not(p91_out);
    p91 : perceptron
        Generic map (
            WEIGHTS => "0000000000000000000000000111111110001111000001100000001000011111111100111000000000100111111111111111111111011111111111",
            SHIFT => 4,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p91_in,
            y(0) => p91_out,
            y(1 to 17 - 1) => dummy91
        );


    p92_in <= x(37) & x(62) & x(63) & x(64) & x(90) & x(108) & x(164) & x(165) & x(166) & x(171) & x(191) & x(192) & x(193) & x(194) & x(199) & x(210) & x(211) & x(218) & x(219) & x(220) & x(221) & x(222) & x(237) & x(238) & x(239) & x(247) & x(248) & x(249) & x(250) & x(266) & x(267) & x(275) & x(276) & x(277) & x(294) & x(295) & x(296) & x(305) & x(306) & x(320) & x(322) & x(323) & x(327) & x(328) & x(330) & x(331) & x(332) & x(347) & x(348) & x(350) & x(361) & x(366) & x(375) & x(376) & x(418) & x(535) & x(611) & x(677) & x(695) & x(706) & x(709) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(736) & x(737) & x(738) & x(739) & x(740) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(748) & x(749) & x(750) & x(764) & x(770) & x(773);
    y(92) <= not(p92_out);
    p92 : perceptron
        Generic map (
            WEIGHTS => "000001000100001110000011100001100011100011111110011100110111111111111111111111111111111",
            SHIFT => 4,
            B => 245,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p92_in,
            y(0) => p92_out,
            y(1 to 16 - 1) => dummy92
        );


    p93_in <= x(108) & x(146) & x(188) & x(192) & x(211) & x(215) & x(220) & x(221) & x(222) & x(242) & x(243) & x(248) & x(249) & x(250) & x(270) & x(276) & x(277) & x(278) & x(291) & x(305) & x(306) & x(319) & x(328) & x(329) & x(330) & x(333) & x(334) & x(342) & x(345) & x(357) & x(358) & x(359) & x(360) & x(371) & x(386) & x(415) & x(416) & x(445) & x(446) & x(451) & x(473) & x(474) & x(479) & x(480) & x(486) & x(487) & x(501) & x(502) & x(507) & x(508) & x(509) & x(514) & x(515) & x(528) & x(529) & x(530) & x(535) & x(537) & x(556) & x(557) & x(558) & x(563) & x(565) & x(583) & x(584) & x(591) & x(593) & x(611) & x(612) & x(619) & x(620) & x(624) & x(640) & x(646) & x(647) & x(648) & x(659) & x(660) & x(692) & x(693) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(742) & x(743) & x(744) & x(746) & x(747) & x(748);
    y(93) <= not(p93_out);
    p93 : perceptron
        Generic map (
            WEIGHTS => "011101111111111111011000011000000000011111110011111001111111111111111111111111000000000000000",
            SHIFT => 4,
            B => 503,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p93_in,
            y(0) => p93_out,
            y(1 to 16 - 1) => dummy93
        );


    p94_in <= x(35) & x(40) & x(44) & x(63) & x(68) & x(69) & x(79) & x(165) & x(166) & x(181) & x(184) & x(185) & x(193) & x(194) & x(199) & x(207) & x(208) & x(209) & x(210) & x(211) & x(212) & x(213) & x(221) & x(243) & x(248) & x(249) & x(250) & x(263) & x(271) & x(274) & x(275) & x(276) & x(277) & x(278) & x(294) & x(295) & x(305) & x(320) & x(328) & x(333) & x(334) & x(347) & x(348) & x(350) & x(353) & x(356) & x(369) & x(376) & x(397) & x(415) & x(416) & x(490) & x(529) & x(541) & x(544) & x(545) & x(557) & x(612) & x(675) & x(692) & x(693) & x(694) & x(695) & x(697) & x(706) & x(707) & x(708) & x(709) & x(715) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(746) & x(747) & x(748) & x(777);
    y(94) <= not(p94_out);
    p94 : perceptron
        Generic map (
            WEIGHTS => "11111110000000000000000000000000001100000001000000011011110000010000000000000001",
            SHIFT => 4,
            B => -441,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p94_in,
            y(0) => p94_out,
            y(1 to 16 - 1) => dummy94
        );


    p95_in <= x(35) & x(37) & x(38) & x(39) & x(40) & x(41) & x(42) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(92) & x(95) & x(96) & x(127) & x(158) & x(166) & x(182) & x(183) & x(193) & x(194) & x(198) & x(221) & x(222) & x(248) & x(249) & x(250) & x(276) & x(277) & x(278) & x(297) & x(305) & x(306) & x(309) & x(311) & x(324) & x(325) & x(326) & x(334) & x(362) & x(381) & x(394) & x(399) & x(408) & x(409) & x(411) & x(434) & x(437) & x(444) & x(464) & x(465) & x(489) & x(541) & x(542) & x(543) & x(570) & x(572) & x(611) & x(641) & x(707) & x(710) & x(719) & x(735) & x(736) & x(737) & x(738) & x(739) & x(740) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(765) & x(770) & x(773);
    y(95) <= not(p95_out);
    p95 : perceptron
        Generic map (
            WEIGHTS => "11111111111111111111111101111111101100000110000001010011111111000000000000000000",
            SHIFT => 4,
            B => 260,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p95_in,
            y(0) => p95_out,
            y(1 to 16 - 1) => dummy95
        );


    p96_in <= x(34) & x(35) & x(37) & x(38) & x(39) & x(40) & x(41) & x(63) & x(64) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(105) & x(106) & x(107) & x(108) & x(135) & x(154) & x(162) & x(163) & x(164) & x(165) & x(192) & x(193) & x(194) & x(195) & x(221) & x(222) & x(248) & x(249) & x(250) & x(277) & x(278) & x(289) & x(290) & x(292) & x(295) & x(302) & x(303) & x(305) & x(312) & x(320) & x(328) & x(329) & x(330) & x(331) & x(332) & x(339) & x(345) & x(353) & x(354) & x(356) & x(357) & x(358) & x(359) & x(360) & x(366) & x(386) & x(387) & x(388) & x(414) & x(418) & x(446) & x(451) & x(473) & x(474) & x(479) & x(485) & x(486) & x(487) & x(497) & x(500) & x(501) & x(502) & x(507) & x(509) & x(513) & x(514) & x(515) & x(525) & x(528) & x(529) & x(530) & x(535) & x(551) & x(556) & x(557) & x(558) & x(563) & x(565) & x(566) & x(580) & x(584) & x(585) & x(591) & x(597) & x(612) & x(613) & x(619) & x(620) & x(624) & x(625) & x(638) & x(640) & x(648) & x(649) & x(657) & x(676) & x(677) & x(678) & x(690) & x(691) & x(692) & x(693) & x(695) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(746) & x(747) & x(748) & x(749) & x(764) & x(765) & x(769) & x(773) & x(774);
    y(96) <= not(p96_out);
    p96 : perceptron
        Generic map (
            WEIGHTS => "111111111111111111110000000000000000011101100111111011111111011110000001110000001110000000000000000000000000001000111111111111111100000",
            SHIFT => 4,
            B => -176,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p96_in,
            y(0) => p96_out,
            y(1 to 17 - 1) => dummy96
        );


    p97_in <= x(34) & x(35) & x(36) & x(37) & x(39) & x(40) & x(41) & x(43) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(79) & x(103) & x(104) & x(105) & x(106) & x(107) & x(108) & x(118) & x(121) & x(151) & x(174) & x(176) & x(195) & x(215) & x(221) & x(222) & x(242) & x(249) & x(250) & x(277) & x(278) & x(283) & x(288) & x(294) & x(295) & x(296) & x(305) & x(311) & x(312) & x(317) & x(319) & x(320) & x(329) & x(330) & x(331) & x(332) & x(338) & x(339) & x(348) & x(357) & x(358) & x(359) & x(360) & x(362) & x(366) & x(380) & x(385) & x(386) & x(387) & x(388) & x(390) & x(403) & x(408) & x(414) & x(415) & x(418) & x(431) & x(444) & x(446) & x(466) & x(473) & x(474) & x(479) & x(485) & x(486) & x(487) & x(500) & x(501) & x(502) & x(507) & x(510) & x(513) & x(514) & x(515) & x(527) & x(528) & x(529) & x(530) & x(535) & x(536) & x(537) & x(551) & x(552) & x(553) & x(555) & x(556) & x(557) & x(558) & x(563) & x(564) & x(566) & x(579) & x(583) & x(584) & x(585) & x(586) & x(591) & x(596) & x(597) & x(610) & x(611) & x(612) & x(613) & x(619) & x(620) & x(625) & x(638) & x(639) & x(640) & x(648) & x(649) & x(650) & x(651) & x(677) & x(688) & x(690) & x(691) & x(692) & x(693) & x(694) & x(695) & x(719) & x(720) & x(721) & x(722) & x(723) & x(750) & x(764) & x(765) & x(766) & x(769) & x(770) & x(773) & x(774);
    y(97) <= not(p97_out);
    p97 : perceptron
        Generic map (
            WEIGHTS => "111111111111111111111111111111110000000000000001000000111111100111110011111011110110000011100000111000000000000000000000000000000000000000011111111111100000000",
            SHIFT => 4,
            B => -190,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p97_in,
            y(0) => p97_out,
            y(1 to 17 - 1) => dummy97
        );


    p98_in <= x(35) & x(40) & x(41) & x(43) & x(66) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(102) & x(103) & x(104) & x(105) & x(106) & x(107) & x(118) & x(121) & x(151) & x(178) & x(181) & x(215) & x(241) & x(267) & x(277) & x(287) & x(290) & x(295) & x(303) & x(318) & x(320) & x(330) & x(331) & x(343) & x(344) & x(348) & x(349) & x(354) & x(355) & x(356) & x(357) & x(358) & x(359) & x(381) & x(386) & x(387) & x(390) & x(406) & x(407) & x(408) & x(414) & x(418) & x(434) & x(446) & x(450) & x(473) & x(474) & x(479) & x(487) & x(500) & x(501) & x(502) & x(507) & x(508) & x(509) & x(513) & x(514) & x(515) & x(516) & x(528) & x(529) & x(530) & x(535) & x(536) & x(537) & x(553) & x(556) & x(557) & x(558) & x(563) & x(564) & x(566) & x(579) & x(580) & x(581) & x(583) & x(584) & x(585) & x(591) & x(592) & x(596) & x(611) & x(612) & x(613) & x(619) & x(620) & x(624) & x(625) & x(637) & x(638) & x(639) & x(640) & x(647) & x(648) & x(649) & x(650) & x(690) & x(691) & x(692) & x(695) & x(708) & x(721) & x(722);
    y(98) <= not(p98_out);
    p98 : perceptron
        Generic map (
            WEIGHTS => "00000000000000000000001111111110010000000000000000001000010111110111111000011111111111111111111111111111111111110000100",
            SHIFT => 4,
            B => 181,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p98_in,
            y(0) => p98_out,
            y(1 to 17 - 1) => dummy98
        );


    p99_in <= x(35) & x(41) & x(97) & x(99) & x(100) & x(101) & x(102) & x(103) & x(106) & x(107) & x(108) & x(163) & x(164) & x(165) & x(166) & x(191) & x(192) & x(193) & x(194) & x(198) & x(199) & x(219) & x(220) & x(221) & x(222) & x(226) & x(227) & x(237) & x(247) & x(248) & x(249) & x(250) & x(251) & x(254) & x(255) & x(256) & x(264) & x(265) & x(266) & x(276) & x(277) & x(278) & x(282) & x(283) & x(284) & x(293) & x(294) & x(305) & x(306) & x(309) & x(310) & x(311) & x(312) & x(329) & x(330) & x(331) & x(332) & x(333) & x(334) & x(337) & x(338) & x(339) & x(349) & x(350) & x(351) & x(359) & x(360) & x(366) & x(376) & x(377) & x(378) & x(386) & x(388) & x(406) & x(414) & x(433) & x(434) & x(441) & x(460) & x(461) & x(463) & x(486) & x(490) & x(499) & x(513) & x(543) & x(557) & x(572) & x(573) & x(601) & x(653) & x(693) & x(694) & x(695) & x(706) & x(707) & x(708) & x(711) & x(712) & x(713) & x(714) & x(735) & x(736) & x(737) & x(739) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(748) & x(764) & x(765) & x(766) & x(769) & x(770) & x(771) & x(772) & x(773) & x(774);
    y(99) <= not(p99_out);
    p99 : perceptron
        Generic map (
            WEIGHTS => "1111111111100000000110000111000001111110001111100111111110011100011100011010010001011111110000111111111111111110111111111",
            SHIFT => 4,
            B => 437,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p99_in,
            y(0) => p99_out,
            y(1 to 17 - 1) => dummy99
        );


    p100_in <= x(35) & x(36) & x(37) & x(38) & x(39) & x(40) & x(41) & x(44) & x(45) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(78) & x(79) & x(90) & x(91) & x(92) & x(93) & x(94) & x(95) & x(96) & x(100) & x(101) & x(102) & x(104) & x(105) & x(136) & x(193) & x(198) & x(219) & x(220) & x(247) & x(248) & x(266) & x(275) & x(294) & x(320) & x(348) & x(353) & x(361) & x(362) & x(380) & x(387) & x(394) & x(396) & x(401) & x(404) & x(408) & x(432) & x(436) & x(442) & x(460) & x(469) & x(479) & x(496) & x(497) & x(507) & x(529) & x(535) & x(557) & x(563) & x(564) & x(591) & x(592) & x(602) & x(619) & x(620) & x(647) & x(648) & x(649) & x(657) & x(676) & x(691) & x(692) & x(718) & x(719) & x(720) & x(721) & x(745) & x(746) & x(747) & x(773);
    y(100) <= not(p100_out);
    p100 : perceptron
        Generic map (
            WEIGHTS => "1111111111111111111111111111111111111100000001010000001001000010111111111111111111010000000000",
            SHIFT => 4,
            B => 727,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p100_in,
            y(0) => p100_out,
            y(1 to 16 - 1) => dummy100
        );


    p101_in <= x(34) & x(35) & x(36) & x(37) & x(38) & x(39) & x(40) & x(41) & x(44) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(75) & x(76) & x(90) & x(91) & x(92) & x(93) & x(94) & x(95) & x(96) & x(102) & x(103) & x(146) & x(171) & x(172) & x(173) & x(197) & x(199) & x(200) & x(221) & x(222) & x(227) & x(228) & x(248) & x(249) & x(250) & x(276) & x(277) & x(297) & x(299) & x(300) & x(367) & x(370) & x(396) & x(397) & x(398) & x(406) & x(409) & x(424) & x(425) & x(433) & x(434) & x(437) & x(445) & x(450) & x(462) & x(473) & x(487) & x(506) & x(507) & x(515) & x(516) & x(534) & x(535) & x(542) & x(543) & x(544) & x(563) & x(573) & x(611) & x(618) & x(619) & x(638) & x(640) & x(647) & x(648) & x(675) & x(676) & x(677) & x(678) & x(679) & x(693) & x(694) & x(695) & x(706) & x(708) & x(709) & x(710) & x(713) & x(736) & x(748);
    y(101) <= not(p101_out);
    p101 : perceptron
        Generic map (
            WEIGHTS => "1111111111111111111111111111111000000011001111100010000100011010111001100111011001100000000000000000",
            SHIFT => 4,
            B => 84,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p101_in,
            y(0) => p101_out,
            y(1 to 16 - 1) => dummy101
        );


    p102_in <= x(63) & x(64) & x(79) & x(104) & x(105) & x(106) & x(107) & x(108) & x(135) & x(162) & x(163) & x(164) & x(165) & x(192) & x(193) & x(194) & x(195) & x(211) & x(220) & x(221) & x(222) & x(248) & x(249) & x(250) & x(276) & x(277) & x(301) & x(302) & x(303) & x(305) & x(326) & x(327) & x(328) & x(329) & x(330) & x(331) & x(332) & x(348) & x(356) & x(357) & x(358) & x(359) & x(360) & x(375) & x(376) & x(386) & x(387) & x(388) & x(418) & x(479) & x(484) & x(495) & x(513) & x(514) & x(515) & x(516) & x(522) & x(523) & x(535) & x(550) & x(551) & x(556) & x(563) & x(578) & x(677) & x(692) & x(695) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(745) & x(746) & x(747) & x(748) & x(749) & x(764);
    y(102) <= not(p102_out);
    p102 : perceptron
        Generic map (
            WEIGHTS => "111111110000000001000000001110111111101111100111001011110000000001111111111111110",
            SHIFT => 4,
            B => 183,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p102_in,
            y(0) => p102_out,
            y(1 to 16 - 1) => dummy102
        );


    p103_in <= x(35) & x(36) & x(38) & x(39) & x(40) & x(41) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(74) & x(75) & x(76) & x(77) & x(78) & x(79) & x(90) & x(91) & x(92) & x(93) & x(94) & x(95) & x(96) & x(97) & x(98) & x(99) & x(100) & x(101) & x(102) & x(103) & x(104) & x(105) & x(106) & x(107) & x(108) & x(163) & x(164) & x(165) & x(191) & x(192) & x(193) & x(210) & x(211) & x(212) & x(219) & x(220) & x(221) & x(222) & x(238) & x(239) & x(248) & x(249) & x(250) & x(276) & x(277) & x(302) & x(303) & x(305) & x(327) & x(328) & x(329) & x(330) & x(331) & x(333) & x(334) & x(338) & x(349) & x(357) & x(358) & x(359) & x(366) & x(400) & x(445) & x(450) & x(473) & x(474) & x(487) & x(501) & x(513) & x(514) & x(515) & x(529) & x(542) & x(543) & x(557) & x(709) & x(713) & x(714) & x(715) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(732) & x(736) & x(737) & x(738) & x(739) & x(740) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(748) & x(749) & x(750) & x(773) & x(774);
    y(103) <= not(p103_out);
    p103 : perceptron
        Generic map (
            WEIGHTS => "00000000000000000000000000000000000000000011111100011110011111001000001101000010100000000000000000000000000000000000000000",
            SHIFT => 4,
            B => -1243,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p103_in,
            y(0) => p103_out,
            y(1 to 17 - 1) => dummy103
        );


    p104_in <= x(37) & x(38) & x(39) & x(40) & x(41) & x(45) & x(46) & x(63) & x(64) & x(66) & x(67) & x(68) & x(69) & x(70) & x(72) & x(73) & x(74) & x(75) & x(76) & x(78) & x(79) & x(104) & x(105) & x(146) & x(163) & x(182) & x(191) & x(192) & x(197) & x(198) & x(212) & x(220) & x(221) & x(222) & x(238) & x(248) & x(249) & x(264) & x(277) & x(291) & x(302) & x(303) & x(304) & x(309) & x(326) & x(328) & x(329) & x(330) & x(331) & x(332) & x(338) & x(349) & x(350) & x(357) & x(361) & x(362) & x(366) & x(390) & x(394) & x(400) & x(414) & x(416) & x(418) & x(438) & x(446) & x(450) & x(462) & x(474) & x(475) & x(478) & x(501) & x(502) & x(506) & x(507) & x(513) & x(514) & x(515) & x(529) & x(534) & x(535) & x(540) & x(557) & x(563) & x(591) & x(592) & x(618) & x(619) & x(620) & x(647) & x(648) & x(649) & x(675) & x(676) & x(677) & x(678) & x(679) & x(692) & x(703) & x(712) & x(713) & x(714) & x(715) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(736) & x(737) & x(738) & x(739) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(748) & x(749) & x(750) & x(764) & x(773);
    y(104) <= not(p104_out);
    p104 : perceptron
        Generic map (
            WEIGHTS => "111111111111111111111111101110011101101000000000000110000001110101100100110000110011111111111111010000000000000000000000000000",
            SHIFT => 4,
            B => 125,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p104_in,
            y(0) => p104_out,
            y(1 to 17 - 1) => dummy104
        );


    p105_in <= x(44) & x(51) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(77) & x(91) & x(93) & x(94) & x(95) & x(96) & x(97) & x(98) & x(105) & x(106) & x(108) & x(182) & x(183) & x(191) & x(192) & x(210) & x(211) & x(212) & x(224) & x(238) & x(239) & x(330) & x(331) & x(335) & x(338) & x(363) & x(390) & x(397) & x(398) & x(414) & x(445) & x(446) & x(447) & x(463) & x(473) & x(474) & x(477) & x(501) & x(502) & x(505) & x(529) & x(533) & x(557) & x(695) & x(709) & x(710) & x(711) & x(712) & x(713) & x(714) & x(715) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(732) & x(737) & x(738) & x(739) & x(740) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(748) & x(749) & x(750);
    y(105) <= not(p105_out);
    p105 : perceptron
        Generic map (
            WEIGHTS => "010000000000000000000001100010000101011100110010010100000000000000000000000000000000",
            SHIFT => 5,
            B => -1301,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p105_in,
            y(0) => p105_out,
            y(1 to 17 - 1) => dummy105
        );


    p106_in <= x(34) & x(35) & x(37) & x(39) & x(40) & x(41) & x(66) & x(68) & x(69) & x(74) & x(165) & x(166) & x(192) & x(193) & x(220) & x(221) & x(247) & x(248) & x(249) & x(250) & x(276) & x(277) & x(305) & x(334) & x(359) & x(362) & x(370) & x(386) & x(387) & x(388) & x(390) & x(400) & x(401) & x(413) & x(414) & x(415) & x(416) & x(418) & x(428) & x(429) & x(446) & x(450) & x(473) & x(474) & x(475) & x(500) & x(501) & x(502) & x(528) & x(529) & x(530) & x(538) & x(556) & x(557) & x(558) & x(566) & x(583) & x(584) & x(595) & x(596) & x(597) & x(611) & x(612) & x(624) & x(625) & x(626) & x(640) & x(657) & x(675) & x(676) & x(677) & x(678) & x(744) & x(746) & x(747) & x(748) & x(770) & x(773);
    y(106) <= not(p106_out);
    p106 : perceptron
        Generic map (
            WEIGHTS => "000000000011111111111111010000100000010010111111111111111111111111110000111111",
            SHIFT => 4,
            B => 425,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p106_in,
            y(0) => p106_out,
            y(1 to 16 - 1) => dummy106
        );


    p107_in <= x(37) & x(38) & x(39) & x(40) & x(41) & x(45) & x(46) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(79) & x(103) & x(104) & x(105) & x(106) & x(118) & x(135) & x(154) & x(164) & x(165) & x(171) & x(181) & x(182) & x(183) & x(191) & x(192) & x(193) & x(200) & x(210) & x(211) & x(219) & x(220) & x(221) & x(238) & x(239) & x(247) & x(248) & x(249) & x(267) & x(276) & x(277) & x(291) & x(292) & x(294) & x(295) & x(296) & x(303) & x(304) & x(316) & x(317) & x(319) & x(320) & x(321) & x(323) & x(326) & x(330) & x(331) & x(332) & x(333) & x(343) & x(344) & x(347) & x(349) & x(350) & x(353) & x(354) & x(355) & x(356) & x(357) & x(358) & x(361) & x(371) & x(372) & x(376) & x(378) & x(381) & x(382) & x(390) & x(391) & x(398) & x(399) & x(400) & x(408) & x(418) & x(426) & x(427) & x(428) & x(429) & x(431) & x(436) & x(446) & x(450) & x(455) & x(456) & x(457) & x(458) & x(459) & x(460) & x(463) & x(464) & x(473) & x(474) & x(475) & x(479) & x(483) & x(484) & x(485) & x(486) & x(487) & x(488) & x(490) & x(491) & x(495) & x(501) & x(502) & x(507) & x(514) & x(515) & x(516) & x(529) & x(534) & x(535) & x(557) & x(558) & x(562) & x(563) & x(564) & x(584) & x(591) & x(619) & x(620) & x(623) & x(624) & x(625) & x(626) & x(627) & x(631) & x(632) & x(647) & x(651) & x(652) & x(653) & x(654) & x(655) & x(656) & x(657) & x(658) & x(659) & x(680) & x(681) & x(682) & x(684) & x(704) & x(717) & x(718) & x(719) & x(720) & x(721) & x(723) & x(745) & x(746) & x(747) & x(748) & x(749);
    y(107) <= not(p107_out);
    p107 : perceptron
        Generic map (
            WEIGHTS => "1111111111111111111111111111101011000011100011100111011110000011110010000111001111110110011001111011111100111111110000111111110000111000000000000000000000000000000000100000000000",
            SHIFT => 3,
            B => 28,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p107_in,
            y(0) => p107_out,
            y(1 to 16 - 1) => dummy107
        );


    p108_in <= x(37) & x(64) & x(66) & x(118) & x(155) & x(182) & x(184) & x(186) & x(218) & x(243) & x(245) & x(246) & x(271) & x(273) & x(274) & x(275) & x(296) & x(297) & x(299) & x(300) & x(301) & x(302) & x(305) & x(333) & x(342) & x(343) & x(347) & x(361) & x(369) & x(370) & x(371) & x(390) & x(391) & x(397) & x(400) & x(401) & x(402) & x(416) & x(418) & x(428) & x(429) & x(446) & x(450) & x(473) & x(474) & x(475) & x(479) & x(501) & x(502) & x(507) & x(528) & x(529) & x(530) & x(535) & x(557) & x(558) & x(563) & x(584) & x(591) & x(597) & x(612) & x(619) & x(640) & x(647) & x(656) & x(657) & x(658) & x(659) & x(720) & x(747);
    y(108) <= not(p108_out);
    p108 : perceptron
        Generic map (
            WEIGHTS => "1110000000000000000000001110111001111101100000000000000000000000000000",
            SHIFT => 4,
            B => -483,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p108_in,
            y(0) => p108_out,
            y(1 to 16 - 1) => dummy108
        );


    p109_in <= x(62) & x(78) & x(103) & x(104) & x(105) & x(106) & x(107) & x(151) & x(152) & x(153) & x(154) & x(155) & x(178) & x(190) & x(191) & x(221) & x(249) & x(250) & x(277) & x(319) & x(325) & x(327) & x(329) & x(330) & x(343) & x(346) & x(352) & x(353) & x(355) & x(370) & x(371) & x(378) & x(398) & x(399) & x(400) & x(405) & x(460) & x(486) & x(487) & x(488) & x(513) & x(514) & x(515) & x(516) & x(542) & x(692) & x(693) & x(695) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(742) & x(746) & x(747) & x(748);
    y(109) <= not(p109_out);
    p109 : perceptron
        Generic map (
            WEIGHTS => "1111111111111000000011110011100100011111111111111111111111",
            SHIFT => 4,
            B => 244,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p109_in,
            y(0) => p109_out,
            y(1 to 16 - 1) => dummy109
        );


    p110_in <= x(64) & x(93) & x(145) & x(172) & x(198) & x(221) & x(226) & x(248) & x(249) & x(250) & x(254) & x(276) & x(277) & x(282) & x(302) & x(303) & x(310) & x(311) & x(322) & x(323) & x(327) & x(329) & x(330) & x(331) & x(332) & x(338) & x(339) & x(348) & x(349) & x(350) & x(351) & x(358) & x(359) & x(360) & x(366) & x(376) & x(377) & x(378) & x(379) & x(390) & x(404) & x(405) & x(406) & x(418) & x(432) & x(433) & x(434) & x(450) & x(460) & x(461) & x(473) & x(474) & x(478) & x(484) & x(487) & x(488) & x(500) & x(501) & x(502) & x(506) & x(507) & x(515) & x(528) & x(529) & x(534) & x(535) & x(556) & x(557) & x(584) & x(611) & x(619) & x(638) & x(646) & x(647) & x(648) & x(675) & x(690) & x(691) & x(692) & x(693) & x(694) & x(695) & x(696) & x(707) & x(708) & x(720) & x(722) & x(723) & x(735) & x(736) & x(737) & x(738) & x(739) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(764) & x(765) & x(766) & x(769) & x(770) & x(772) & x(773) & x(774);
    y(110) <= not(p110_out);
    p110 : perceptron
        Generic map (
            WEIGHTS => "11001111111111001100000001100000001000010001000000110000111000110011110100000000000110001111111111111111111",
            SHIFT => 4,
            B => 224,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p110_in,
            y(0) => p110_out,
            y(1 to 16 - 1) => dummy110
        );


    p111_in <= x(37) & x(40) & x(49) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(92) & x(104) & x(105) & x(106) & x(118) & x(124) & x(135) & x(154) & x(164) & x(165) & x(166) & x(171) & x(172) & x(173) & x(174) & x(191) & x(192) & x(193) & x(194) & x(219) & x(220) & x(221) & x(222) & x(247) & x(248) & x(249) & x(250) & x(254) & x(260) & x(263) & x(276) & x(277) & x(278) & x(287) & x(289) & x(290) & x(291) & x(292) & x(295) & x(296) & x(297) & x(298) & x(300) & x(302) & x(305) & x(306) & x(317) & x(319) & x(320) & x(330) & x(331) & x(332) & x(340) & x(341) & x(342) & x(343) & x(344) & x(348) & x(359) & x(360) & x(366) & x(368) & x(394) & x(424) & x(425) & x(428) & x(429) & x(439) & x(440) & x(446) & x(450) & x(453) & x(454) & x(456) & x(474) & x(502) & x(529) & x(534) & x(535) & x(557) & x(558) & x(563) & x(584) & x(591) & x(612) & x(619) & x(642) & x(647) & x(685) & x(706) & x(707) & x(708) & x(709) & x(710) & x(711) & x(712) & x(713) & x(715) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(736) & x(737) & x(738) & x(739) & x(740) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(748) & x(764) & x(765) & x(766) & x(770) & x(773);
    y(111) <= not(p111_out);
    p111 : perceptron
        Generic map (
            WEIGHTS => "11111111111111100101110000111111111111111111111110000001111100011111100111000000000000000000000000011111111111111111111111111111111111",
            SHIFT => 4,
            B => 752,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p111_in,
            y(0) => p111_out,
            y(1 to 17 - 1) => dummy111
        );


    p112_in <= x(40) & x(41) & x(152) & x(155) & x(156) & x(171) & x(178) & x(179) & x(180) & x(181) & x(192) & x(193) & x(207) & x(208) & x(209) & x(219) & x(247) & x(248) & x(290) & x(291) & x(294) & x(295) & x(322) & x(348) & x(360) & x(372) & x(376) & x(400) & x(414) & x(416) & x(432) & x(433) & x(446) & x(450) & x(460) & x(473) & x(486) & x(487) & x(488) & x(500) & x(501) & x(502) & x(506) & x(513) & x(514) & x(515) & x(516) & x(528) & x(529) & x(530) & x(534) & x(535) & x(540) & x(552) & x(556) & x(557) & x(566) & x(567) & x(568) & x(569) & x(583) & x(584) & x(595) & x(596) & x(597) & x(598) & x(607) & x(611) & x(626) & x(627) & x(656) & x(675) & x(676) & x(677) & x(678) & x(679) & x(705) & x(706) & x(708) & x(719) & x(720) & x(721) & x(723);
    y(112) <= not(p112_out);
    p112 : perceptron
        Generic map (
            WEIGHTS => "11000100000000000000111011011100010000000010000000110000000000000000000111111111111",
            SHIFT => 3,
            B => -76,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p112_in,
            y(0) => p112_out,
            y(1 to 15 - 1) => dummy112
        );


    p113_in <= x(35) & x(38) & x(39) & x(44) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(78) & x(79) & x(90) & x(91) & x(92) & x(93) & x(94) & x(95) & x(96) & x(104) & x(105) & x(106) & x(171) & x(172) & x(193) & x(199) & x(200) & x(227) & x(247) & x(248) & x(249) & x(264) & x(267) & x(275) & x(276) & x(277) & x(291) & x(292) & x(294) & x(295) & x(296) & x(306) & x(322) & x(323) & x(324) & x(350) & x(351) & x(370) & x(378) & x(397) & x(425) & x(432) & x(445) & x(450) & x(460) & x(473) & x(474) & x(487) & x(488) & x(500) & x(501) & x(506) & x(507) & x(513) & x(514) & x(515) & x(516) & x(528) & x(529) & x(534) & x(535) & x(541) & x(542) & x(543) & x(556) & x(557) & x(563) & x(583) & x(584) & x(610) & x(611) & x(612) & x(638) & x(640) & x(647) & x(648) & x(675) & x(676) & x(677) & x(678) & x(706) & x(720);
    y(113) <= not(p113_out);
    p113 : perceptron
        Generic map (
            WEIGHTS => "00000000000000000000000001101110000100000111011111111100100000001100000011000001000000011111110",
            SHIFT => 4,
            B => -447,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p113_in,
            y(0) => p113_out,
            y(1 to 16 - 1) => dummy113
        );


    p114_in <= x(104) & x(105) & x(106) & x(107) & x(151) & x(152) & x(177) & x(182) & x(198) & x(210) & x(221) & x(222) & x(248) & x(249) & x(250) & x(276) & x(277) & x(278) & x(305) & x(306) & x(309) & x(310) & x(311) & x(326) & x(329) & x(330) & x(337) & x(338) & x(339) & x(350) & x(357) & x(366) & x(378) & x(450) & x(479) & x(484) & x(485) & x(506) & x(507) & x(514) & x(515) & x(516) & x(535) & x(563) & x(566) & x(591) & x(592) & x(595) & x(596) & x(619) & x(620) & x(623) & x(624) & x(625) & x(647) & x(648) & x(649) & x(655) & x(656) & x(657) & x(658) & x(675) & x(676) & x(677) & x(694) & x(695) & x(719) & x(720) & x(721) & x(723) & x(748) & x(749) & x(769) & x(770) & x(771) & x(773) & x(774);
    y(114) <= not(p114_out);
    p114 : perceptron
        Generic map (
            WEIGHTS => "00001111011111111111000000000100111001100011111111111111111111111111111100000",
            SHIFT => 4,
            B => 316,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p114_in,
            y(0) => p114_out,
            y(1 to 16 - 1) => dummy114
        );


    p115_in <= x(14) & x(71) & x(72) & x(73) & x(79) & x(81) & x(86) & x(114) & x(252) & x(283) & x(295) & x(303) & x(321) & x(322) & x(331) & x(333) & x(334) & x(339) & x(348) & x(349) & x(350) & x(351) & x(361) & x(365) & x(366) & x(376) & x(377) & x(378) & x(379) & x(393) & x(405) & x(406) & x(433) & x(473) & x(501) & x(502) & x(528) & x(529) & x(556) & x(557) & x(584) & x(586) & x(611) & x(612) & x(638) & x(642) & x(656) & x(657) & x(674) & x(691) & x(692) & x(693) & x(694) & x(695) & x(708) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(736) & x(748) & x(764) & x(766) & x(770) & x(771) & x(773) & x(774);
    y(115) <= not(p115_out);
    p115 : perceptron
        Generic map (
            WEIGHTS => "100011111110000001000001100001000111111111111100100000100000010111111",
            SHIFT => 4,
            B => -720,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p115_in,
            y(0) => p115_out,
            y(1 to 16 - 1) => dummy115
        );


    p116_in <= x(35) & x(36) & x(37) & x(38) & x(39) & x(40) & x(41) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(78) & x(90) & x(91) & x(92) & x(93) & x(97) & x(105) & x(106) & x(127) & x(145) & x(146) & x(171) & x(172) & x(173) & x(174) & x(182) & x(197) & x(199) & x(200) & x(201) & x(202) & x(205) & x(210) & x(211) & x(212) & x(227) & x(228) & x(229) & x(231) & x(232) & x(249) & x(250) & x(256) & x(276) & x(277) & x(297) & x(299) & x(311) & x(312) & x(324) & x(333) & x(348) & x(353) & x(358) & x(361) & x(376) & x(381) & x(386) & x(387) & x(422) & x(423) & x(436) & x(450) & x(464) & x(465) & x(475) & x(478) & x(479) & x(492) & x(506) & x(507) & x(514) & x(515) & x(534) & x(535) & x(539) & x(542) & x(563) & x(570) & x(591) & x(618) & x(619) & x(647) & x(648) & x(657) & x(675) & x(676) & x(677) & x(681) & x(682) & x(683) & x(684) & x(692) & x(693) & x(694) & x(695) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(732) & x(742) & x(746) & x(747) & x(748) & x(749) & x(769) & x(770) & x(771) & x(773);
    y(116) <= not(p116_out);
    p116 : perceptron
        Generic map (
            WEIGHTS => "00000000000000000000000000011111101111110001111100100111111110111001111111111110011001011111111111110000000000000000001111",
            SHIFT => 4,
            B => -98,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p116_in,
            y(0) => p116_out,
            y(1 to 17 - 1) => dummy116
        );


    p117_in <= x(0) & x(1) & x(5) & x(7) & x(17) & x(25) & x(26) & x(30) & x(32) & x(33) & x(52) & x(54) & x(55) & x(56) & x(58) & x(59) & x(75) & x(82) & x(105) & x(113) & x(139) & x(141) & x(161) & x(162) & x(165) & x(189) & x(193) & x(198) & x(199) & x(200) & x(201) & x(203) & x(207) & x(217) & x(221) & x(226) & x(227) & x(228) & x(232) & x(233) & x(235) & x(236) & x(242) & x(243) & x(244) & x(249) & x(250) & x(254) & x(255) & x(256) & x(258) & x(267) & x(269) & x(271) & x(276) & x(277) & x(278) & x(282) & x(283) & x(284) & x(293) & x(295) & x(296) & x(309) & x(310) & x(311) & x(312) & x(321) & x(338) & x(339) & x(348) & x(350) & x(355) & x(362) & x(366) & x(367) & x(378) & x(379) & x(382) & x(383) & x(390) & x(405) & x(406) & x(415) & x(418) & x(429) & x(432) & x(433) & x(434) & x(435) & x(459) & x(460) & x(461) & x(462) & x(463) & x(467) & x(468) & x(476) & x(484) & x(486) & x(487) & x(488) & x(489) & x(490) & x(495) & x(503) & x(513) & x(514) & x(515) & x(516) & x(518) & x(529) & x(532) & x(535) & x(546) & x(557) & x(560) & x(584) & x(587) & x(588) & x(611) & x(612) & x(615) & x(616) & x(617) & x(624) & x(643) & x(644) & x(645) & x(651) & x(654) & x(656) & x(657) & x(673) & x(675) & x(676) & x(677) & x(678) & x(679) & x(680) & x(681) & x(690) & x(692) & x(693) & x(694) & x(695) & x(696) & x(704) & x(705) & x(706) & x(707) & x(708) & x(709) & x(710) & x(711) & x(719) & x(720) & x(721) & x(722) & x(723) & x(727) & x(730) & x(735) & x(736) & x(737) & x(743) & x(744) & x(748) & x(749) & x(760) & x(764) & x(765) & x(766) & x(769) & x(770) & x(771) & x(772) & x(773) & x(774) & x(780) & x(781);
    y(117) <= not(p117_out);
    p117 : perceptron
        Generic map (
            WEIGHTS => "1111111111111111111111000000000000000000000000000000000000000000000000011000111101100111111111100111111101111111101111111111101110000100000001111110000000011111110000011100000000011",
            SHIFT => 3,
            B => -63,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p117_in,
            y(0) => p117_out,
            y(1 to 16 - 1) => dummy117
        );


    p118_in <= x(0) & x(1) & x(2) & x(3) & x(4) & x(5) & x(6) & x(7) & x(8) & x(9) & x(10) & x(11) & x(12) & x(15) & x(16) & x(17) & x(18) & x(19) & x(20) & x(21) & x(22) & x(23) & x(24) & x(25) & x(26) & x(27) & x(28) & x(29) & x(30) & x(31) & x(32) & x(33) & x(52) & x(53) & x(54) & x(55) & x(56) & x(57) & x(58) & x(59) & x(61) & x(72) & x(73) & x(74) & x(75) & x(76) & x(82) & x(83) & x(84) & x(85) & x(87) & x(88) & x(104) & x(110) & x(111) & x(112) & x(113) & x(115) & x(136) & x(139) & x(140) & x(141) & x(142) & x(164) & x(165) & x(166) & x(167) & x(168) & x(169) & x(191) & x(192) & x(193) & x(194) & x(196) & x(197) & x(199) & x(219) & x(220) & x(221) & x(222) & x(227) & x(247) & x(248) & x(249) & x(250) & x(251) & x(274) & x(275) & x(276) & x(277) & x(278) & x(304) & x(305) & x(306) & x(307) & x(320) & x(321) & x(322) & x(333) & x(334) & x(347) & x(348) & x(349) & x(350) & x(351) & x(358) & x(359) & x(360) & x(361) & x(362) & x(364) & x(376) & x(377) & x(387) & x(389) & x(392) & x(394) & x(400) & x(401) & x(419) & x(420) & x(427) & x(428) & x(429) & x(448) & x(449) & x(450) & x(451) & x(455) & x(456) & x(476) & x(478) & x(479) & x(501) & x(502) & x(503) & x(504) & x(506) & x(507) & x(529) & x(532) & x(534) & x(535) & x(557) & x(560) & x(563) & x(587) & x(588) & x(591) & x(615) & x(616) & x(617) & x(643) & x(644) & x(645) & x(666) & x(671) & x(672) & x(673) & x(675) & x(677) & x(679) & x(697) & x(698) & x(699) & x(700) & x(701) & x(702) & x(706) & x(707) & x(725) & x(726) & x(727) & x(728) & x(729) & x(730) & x(731) & x(752) & x(753) & x(754) & x(755) & x(756) & x(757) & x(758) & x(759) & x(760) & x(765) & x(770) & x(771) & x(772) & x(773) & x(779) & x(780) & x(781) & x(782) & x(783);
    y(118) <= not(p118_out);
    p118 : perceptron
        Generic map (
            WEIGHTS => "1111111111111111111111111111111111111111100000111111011111011110001110000100000000000000000000000000000001110010010101111111110011100111100110011011011111111110001111110011111111111111110000011111",
            SHIFT => 4,
            B => 946,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p118_in,
            y(0) => p118_out,
            y(1 to 17 - 1) => dummy118
        );


    p119_in <= x(35) & x(37) & x(38) & x(39) & x(40) & x(41) & x(45) & x(46) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(79) & x(101) & x(102) & x(103) & x(104) & x(105) & x(106) & x(192) & x(198) & x(208) & x(212) & x(237) & x(240) & x(263) & x(269) & x(277) & x(291) & x(298) & x(302) & x(303) & x(305) & x(306) & x(329) & x(350) & x(366) & x(378) & x(390) & x(406) & x(418) & x(427) & x(434) & x(439) & x(446) & x(450) & x(451) & x(461) & x(462) & x(474) & x(479) & x(489) & x(490) & x(501) & x(502) & x(507) & x(530) & x(535) & x(557) & x(591) & x(647) & x(648) & x(675) & x(707) & x(709) & x(710) & x(711) & x(712) & x(713) & x(714) & x(715) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(735) & x(736) & x(737) & x(738) & x(739) & x(740) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(769) & x(773);
    y(119) <= not(p119_out);
    p119 : perceptron
        Generic map (
            WEIGHTS => "111111111111111111111111111111111000000010000110101010111011110111001010111100000000000000000000000000000",
            SHIFT => 4,
            B => 109,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p119_in,
            y(0) => p119_out,
            y(1 to 16 - 1) => dummy119
        );


    p120_in <= x(91) & x(93) & x(108) & x(246) & x(294) & x(295) & x(305) & x(306) & x(405) & x(406) & x(416) & x(432) & x(433) & x(450) & x(460) & x(461) & x(473) & x(487) & x(488) & x(489) & x(501) & x(506) & x(514) & x(515) & x(516) & x(528) & x(529) & x(530) & x(557) & x(558) & x(583) & x(584) & x(611) & x(612) & x(626) & x(627) & x(656) & x(657) & x(658) & x(659) & x(675) & x(676) & x(677) & x(678) & x(705) & x(706) & x(719) & x(720) & x(721);
    y(120) <= not(p120_out);
    p120 : perceptron
        Generic map (
            WEIGHTS => "0010110000100100000001000000000000000000111111111",
            SHIFT => 4,
            B => -99,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p120_in,
            y(0) => p120_out,
            y(1 to 15 - 1) => dummy120
        );


    p121_in <= x(66) & x(91) & x(92) & x(93) & x(94) & x(108) & x(145) & x(171) & x(172) & x(173) & x(174) & x(199) & x(200) & x(201) & x(202) & x(227) & x(228) & x(247) & x(248) & x(249) & x(250) & x(255) & x(256) & x(267) & x(276) & x(277) & x(283) & x(284) & x(291) & x(294) & x(295) & x(296) & x(297) & x(299) & x(302) & x(306) & x(309) & x(310) & x(311) & x(322) & x(323) & x(332) & x(337) & x(338) & x(339) & x(357) & x(358) & x(361) & x(362) & x(366) & x(385) & x(387) & x(403) & x(422) & x(450) & x(458) & x(460) & x(478) & x(479) & x(484) & x(485) & x(486) & x(506) & x(507) & x(513) & x(514) & x(515) & x(534) & x(535) & x(543) & x(562) & x(563) & x(591) & x(611) & x(618) & x(619) & x(647) & x(648) & x(650) & x(665) & x(666) & x(675) & x(676) & x(677) & x(678) & x(679) & x(692) & x(706) & x(707) & x(721) & x(732) & x(764) & x(765) & x(769) & x(770) & x(771) & x(772) & x(773) & x(774);
    y(121) <= not(p121_out);
    p121 : perceptron
        Generic map (
            WEIGHTS => "111110000000000001111000110010000001000000000110001110011001110011100100010000011000001001100000000",
            SHIFT => 4,
            B => -549,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p121_in,
            y(0) => p121_out,
            y(1 to 16 - 1) => dummy121
        );


    p122_in <= x(34) & x(35) & x(37) & x(39) & x(40) & x(43) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(71) & x(72) & x(75) & x(103) & x(118) & x(123) & x(124) & x(151) & x(161) & x(164) & x(165) & x(166) & x(171) & x(172) & x(173) & x(174) & x(176) & x(177) & x(192) & x(193) & x(194) & x(197) & x(199) & x(200) & x(201) & x(208) & x(213) & x(220) & x(221) & x(222) & x(228) & x(235) & x(248) & x(249) & x(250) & x(267) & x(269) & x(276) & x(277) & x(296) & x(297) & x(298) & x(299) & x(300) & x(301) & x(302) & x(305) & x(306) & x(311) & x(316) & x(317) & x(318) & x(327) & x(329) & x(331) & x(332) & x(342) & x(343) & x(344) & x(349) & x(350) & x(360) & x(366) & x(370) & x(378) & x(390) & x(405) & x(406) & x(425) & x(434) & x(446) & x(450) & x(453) & x(459) & x(462) & x(473) & x(474) & x(493) & x(501) & x(502) & x(507) & x(528) & x(529) & x(530) & x(534) & x(535) & x(543) & x(556) & x(557) & x(558) & x(562) & x(563) & x(564) & x(565) & x(566) & x(580) & x(584) & x(591) & x(592) & x(612) & x(618) & x(619) & x(620) & x(622) & x(647) & x(675) & x(676) & x(677) & x(691) & x(692) & x(693) & x(694) & x(695) & x(713) & x(719) & x(720) & x(721) & x(722) & x(723) & x(774);
    y(122) <= not(p122_out);
    p122 : perceptron
        Generic map (
            WEIGHTS => "11111111111111111100001111000000111000000111001110011000000011011100001111100110110100011000000000001000000000000000000000111110111110",
            SHIFT => 4,
            B => -155,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p122_in,
            y(0) => p122_out,
            y(1 to 17 - 1) => dummy122
        );


    p123_in <= x(37) & x(38) & x(39) & x(40) & x(41) & x(46) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(79) & x(102) & x(103) & x(104) & x(105) & x(106) & x(157) & x(198) & x(226) & x(227) & x(254) & x(255) & x(256) & x(257) & x(266) & x(267) & x(270) & x(280) & x(282) & x(283) & x(284) & x(285) & x(294) & x(295) & x(305) & x(307) & x(309) & x(310) & x(311) & x(312) & x(319) & x(320) & x(338) & x(339) & x(347) & x(361) & x(362) & x(366) & x(367) & x(376) & x(377) & x(381) & x(382) & x(389) & x(390) & x(394) & x(401) & x(403) & x(404) & x(409) & x(418) & x(430) & x(431) & x(436) & x(446) & x(474) & x(482) & x(502) & x(598) & x(675) & x(693) & x(694) & x(695) & x(696) & x(719) & x(720) & x(721) & x(722) & x(723) & x(735) & x(743) & x(748) & x(749) & x(761) & x(764) & x(765) & x(766) & x(769) & x(770) & x(771) & x(772) & x(773) & x(774);
    y(123) <= not(p123_out);
    p123 : perceptron
        Generic map (
            WEIGHTS => "000000000000000000000000000011111111111111111101111100110111100001110000100011111000000000011001111111111",
            SHIFT => 4,
            B => -8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p123_in,
            y(0) => p123_out,
            y(1 to 16 - 1) => dummy123
        );


    p124_in <= x(108) & x(163) & x(182) & x(183) & x(192) & x(210) & x(211) & x(212) & x(238) & x(239) & x(240) & x(303) & x(315) & x(329) & x(330) & x(331) & x(350) & x(356) & x(357) & x(358) & x(359) & x(416) & x(446) & x(450) & x(487) & x(514) & x(515) & x(535) & x(556) & x(584) & x(677) & x(689) & x(690) & x(691) & x(692) & x(695) & x(715) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(740) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(748) & x(749);
    y(124) <= not(p124_out);
    p124 : perceptron
        Generic map (
            WEIGHTS => "1011011111111111111110101110000111111111111111111111111",
            SHIFT => 4,
            B => 559,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p124_in,
            y(0) => p124_out,
            y(1 to 15 - 1) => dummy124
        );


    p125_in <= x(0) & x(2) & x(12) & x(20) & x(21) & x(33) & x(37) & x(38) & x(39) & x(40) & x(44) & x(45) & x(49) & x(54) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(87) & x(88) & x(112) & x(163) & x(165) & x(177) & x(188) & x(192) & x(194) & x(198) & x(221) & x(222) & x(248) & x(249) & x(250) & x(265) & x(276) & x(277) & x(278) & x(289) & x(291) & x(292) & x(299) & x(301) & x(302) & x(303) & x(305) & x(317) & x(326) & x(327) & x(328) & x(329) & x(330) & x(331) & x(332) & x(350) & x(356) & x(357) & x(358) & x(359) & x(360) & x(378) & x(399) & x(400) & x(419) & x(428) & x(446) & x(450) & x(479) & x(484) & x(485) & x(487) & x(507) & x(513) & x(514) & x(515) & x(532) & x(534) & x(535) & x(563) & x(564) & x(591) & x(592) & x(596) & x(616) & x(617) & x(619) & x(620) & x(624) & x(625) & x(648) & x(649) & x(675) & x(676) & x(677) & x(678) & x(690) & x(691) & x(700) & x(703) & x(705) & x(713) & x(714) & x(715) & x(716) & x(737) & x(738) & x(739) & x(740) & x(741) & x(742) & x(743) & x(752) & x(757) & x(758) & x(759) & x(781);
    y(125) <= not(p125_out);
    p125 : perceptron
        Generic map (
            WEIGHTS => "000000111111101111111110001111110111110111000000010000000010000011101011000100001111111001111111111000110000000000000000",
            SHIFT => 4,
            B => 58,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p125_in,
            y(0) => p125_out,
            y(1 to 17 - 1) => dummy125
        );


    p126_in <= x(34) & x(35) & x(37) & x(38) & x(39) & x(40) & x(41) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(78) & x(79) & x(90) & x(91) & x(93) & x(95) & x(96) & x(97) & x(100) & x(105) & x(129) & x(136) & x(153) & x(165) & x(166) & x(192) & x(193) & x(194) & x(220) & x(221) & x(235) & x(245) & x(247) & x(248) & x(249) & x(250) & x(260) & x(262) & x(263) & x(269) & x(276) & x(277) & x(278) & x(287) & x(290) & x(291) & x(295) & x(305) & x(306) & x(307) & x(313) & x(314) & x(315) & x(316) & x(317) & x(318) & x(319) & x(333) & x(334) & x(340) & x(347) & x(348) & x(350) & x(359) & x(362) & x(368) & x(376) & x(378) & x(387) & x(394) & x(418) & x(440) & x(446) & x(489) & x(523) & x(525) & x(529) & x(535) & x(543) & x(544) & x(545) & x(549) & x(550) & x(552) & x(553) & x(557) & x(563) & x(564) & x(574) & x(576) & x(584) & x(591) & x(612) & x(619) & x(620) & x(648) & x(650) & x(693) & x(697) & x(706) & x(707) & x(708) & x(709) & x(712) & x(713) & x(718) & x(719) & x(720) & x(721) & x(722) & x(735) & x(736) & x(737) & x(739) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(748) & x(750) & x(764) & x(770) & x(773);
    y(126) <= not(p126_out);
    p126 : perceptron
        Generic map (
            WEIGHTS => "111111111111111111111111111111101000000000000000000000001000000000000000110001100101111111111111111111111110100000000000000000000000000",
            SHIFT => 4,
            B => -114,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p126_in,
            y(0) => p126_out,
            y(1 to 17 - 1) => dummy126
        );


    p127_in <= x(44) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(70) & x(91) & x(92) & x(93) & x(94) & x(95) & x(96) & x(135) & x(136) & x(163) & x(171) & x(192) & x(195) & x(199) & x(227) & x(228) & x(294) & x(305) & x(321) & x(322) & x(323) & x(324) & x(333) & x(349) & x(352) & x(361) & x(366) & x(409) & x(423) & x(472) & x(473) & x(474) & x(500) & x(501) & x(502) & x(514) & x(515) & x(528) & x(529) & x(535) & x(541) & x(542) & x(543) & x(556) & x(557) & x(584) & x(611) & x(612) & x(638) & x(675) & x(676) & x(677) & x(678) & x(679) & x(706) & x(707) & x(708) & x(764) & x(770) & x(773);
    y(127) <= not(p127_out);
    p127 : perceptron
        Generic map (
            WEIGHTS => "0000000000000011111111111111111111110000000000100000000011111111111",
            SHIFT => 4,
            B => -57,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p127_in,
            y(0) => p127_out,
            y(1 to 16 - 1) => dummy127
        );


    p128_in <= x(79) & x(108) & x(135) & x(164) & x(165) & x(166) & x(191) & x(192) & x(193) & x(194) & x(219) & x(220) & x(221) & x(222) & x(247) & x(248) & x(249) & x(250) & x(266) & x(267) & x(276) & x(277) & x(278) & x(294) & x(295) & x(297) & x(298) & x(300) & x(301) & x(302) & x(303) & x(305) & x(306) & x(309) & x(328) & x(329) & x(330) & x(331) & x(332) & x(333) & x(334) & x(337) & x(338) & x(348) & x(349) & x(350) & x(357) & x(358) & x(359) & x(360) & x(366) & x(375) & x(376) & x(377) & x(378) & x(381) & x(388) & x(404) & x(405) & x(406) & x(409) & x(436) & x(437) & x(451) & x(474) & x(501) & x(502) & x(514) & x(518) & x(529) & x(545) & x(557) & x(558) & x(584) & x(716) & x(732) & x(744) & x(745) & x(746) & x(773) & x(774);
    y(128) <= not(p128_out);
    p128 : perceptron
        Generic map (
            WEIGHTS => "001111111111111111001110000000011000000110011100000111110111111100000000000000000",
            SHIFT => 4,
            B => -97,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p128_in,
            y(0) => p128_out,
            y(1 to 16 - 1) => dummy128
        );


    p129_in <= x(78) & x(96) & x(97) & x(102) & x(103) & x(105) & x(106) & x(107) & x(108) & x(164) & x(165) & x(166) & x(191) & x(192) & x(193) & x(194) & x(198) & x(219) & x(220) & x(221) & x(222) & x(224) & x(247) & x(248) & x(249) & x(250) & x(251) & x(266) & x(267) & x(276) & x(277) & x(278) & x(297) & x(298) & x(302) & x(305) & x(306) & x(309) & x(310) & x(327) & x(328) & x(329) & x(330) & x(331) & x(332) & x(333) & x(334) & x(338) & x(348) & x(349) & x(350) & x(351) & x(357) & x(359) & x(360) & x(366) & x(377) & x(378) & x(405) & x(406) & x(433) & x(474) & x(500) & x(501) & x(502) & x(514) & x(515) & x(528) & x(529) & x(544) & x(557) & x(584) & x(612) & x(655) & x(681) & x(706) & x(708) & x(716) & x(717) & x(719) & x(732) & x(735) & x(736) & x(737) & x(738) & x(739) & x(740) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(764) & x(766) & x(770) & x(772) & x(773) & x(774);
    y(129) <= not(p129_out);
    p129 : perceptron
        Generic map (
            WEIGHTS => "0000000001111111011111111110011100011000000001101111000011111000000000000110000000000000000000000000",
            SHIFT => 4,
            B => -486,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p129_in,
            y(0) => p129_out,
            y(1 to 16 - 1) => dummy129
        );


    p130_in <= x(35) & x(36) & x(37) & x(38) & x(39) & x(40) & x(41) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(79) & x(90) & x(91) & x(97) & x(100) & x(101) & x(102) & x(103) & x(104) & x(105) & x(106) & x(107) & x(108) & x(136) & x(163) & x(164) & x(165) & x(166) & x(180) & x(191) & x(192) & x(193) & x(194) & x(207) & x(218) & x(219) & x(220) & x(221) & x(222) & x(246) & x(247) & x(248) & x(249) & x(250) & x(274) & x(275) & x(276) & x(277) & x(294) & x(295) & x(303) & x(305) & x(307) & x(320) & x(333) & x(334) & x(347) & x(348) & x(349) & x(358) & x(359) & x(361) & x(362) & x(376) & x(387) & x(390) & x(418) & x(446) & x(490) & x(518) & x(543) & x(544) & x(551) & x(579) & x(656) & x(657) & x(658) & x(719) & x(720) & x(721);
    y(130) <= not(p130_out);
    p130 : perceptron
        Generic map (
            WEIGHTS => "0000000000000000000000000000000000000111111111111111111111111100111111111001110111000011111000",
            SHIFT => 4,
            B => -126,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p130_in,
            y(0) => p130_out,
            y(1 to 16 - 1) => dummy130
        );


    p131_in <= x(37) & x(39) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(70) & x(78) & x(79) & x(91) & x(94) & x(95) & x(96) & x(100) & x(105) & x(106) & x(126) & x(146) & x(147) & x(150) & x(151) & x(174) & x(202) & x(220) & x(247) & x(248) & x(249) & x(277) & x(288) & x(294) & x(305) & x(322) & x(323) & x(333) & x(334) & x(349) & x(350) & x(357) & x(358) & x(360) & x(361) & x(362) & x(387) & x(388) & x(428) & x(429) & x(430) & x(455) & x(456) & x(472) & x(473) & x(501) & x(529) & x(549) & x(557) & x(657) & x(721) & x(748);
    y(131) <= not(p131_out);
    p131 : perceptron
        Generic map (
            WEIGHTS => "000000000000000000000000011111111111111000110000000000000100",
            SHIFT => 4,
            B => -433,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p131_in,
            y(0) => p131_out,
            y(1 to 16 - 1) => dummy131
        );


    p132_in <= x(34) & x(35) & x(37) & x(38) & x(39) & x(40) & x(41) & x(43) & x(44) & x(45) & x(62) & x(63) & x(64) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(79) & x(95) & x(96) & x(97) & x(98) & x(99) & x(100) & x(101) & x(102) & x(103) & x(104) & x(105) & x(106) & x(107) & x(108) & x(162) & x(197) & x(207) & x(242) & x(269) & x(270) & x(284) & x(295) & x(321) & x(323) & x(350) & x(378) & x(386) & x(387) & x(403) & x(414) & x(418) & x(431) & x(446) & x(450) & x(458) & x(515) & x(542) & x(543) & x(548) & x(575) & x(709) & x(710) & x(711) & x(737) & x(738) & x(739) & x(740) & x(741) & x(742) & x(743) & x(744) & x(745);
    y(132) <= not(p132_out);
    p132 : perceptron
        Generic map (
            WEIGHTS => "0000000000000000000000000000000000000000010011101011100001010000000000000000000",
            SHIFT => 4,
            B => -997,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p132_in,
            y(0) => p132_out,
            y(1 to 16 - 1) => dummy132
        );


    p133_in <= x(108) & x(118) & x(133) & x(134) & x(135) & x(154) & x(155) & x(185) & x(197) & x(198) & x(207) & x(217) & x(226) & x(248) & x(249) & x(275) & x(303) & x(304) & x(322) & x(323) & x(329) & x(330) & x(331) & x(332) & x(334) & x(342) & x(350) & x(351) & x(360) & x(361) & x(362) & x(368) & x(370) & x(378) & x(382) & x(390) & x(394) & x(409) & x(410) & x(411) & x(450) & x(474) & x(507) & x(509) & x(526) & x(534) & x(535) & x(539) & x(540) & x(541) & x(542) & x(554) & x(555) & x(557) & x(563) & x(566) & x(567) & x(568) & x(581) & x(582) & x(591) & x(594) & x(598) & x(607) & x(608) & x(610) & x(618) & x(619) & x(646) & x(647) & x(656) & x(674) & x(675) & x(706) & x(708) & x(709) & x(710) & x(711) & x(712) & x(718) & x(719) & x(721) & x(722) & x(735) & x(736) & x(737) & x(738) & x(739) & x(740) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(764) & x(769) & x(770) & x(773);
    y(133) <= not(p133_out);
    p133 : perceptron
        Generic map (
            WEIGHTS => "110001111011011111001111100011100001000011111111111111111111111111111111100000000000000000000000000",
            SHIFT => 4,
            B => 137,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p133_in,
            y(0) => p133_out,
            y(1 to 16 - 1) => dummy133
        );


    p134_in <= x(35) & x(37) & x(38) & x(39) & x(40) & x(41) & x(44) & x(45) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(79) & x(90) & x(91) & x(92) & x(93) & x(94) & x(95) & x(96) & x(100) & x(101) & x(102) & x(103) & x(104) & x(105) & x(106) & x(151) & x(154) & x(181) & x(221) & x(222) & x(248) & x(249) & x(250) & x(276) & x(277) & x(278) & x(289) & x(291) & x(298) & x(299) & x(301) & x(302) & x(305) & x(306) & x(318) & x(322) & x(329) & x(330) & x(332) & x(342) & x(344) & x(345) & x(350) & x(369) & x(373) & x(378) & x(396) & x(397) & x(418) & x(423) & x(425) & x(433) & x(434) & x(445) & x(450) & x(451) & x(473) & x(479) & x(497) & x(507) & x(523) & x(526) & x(535) & x(542) & x(543) & x(550) & x(552) & x(563) & x(584) & x(591) & x(619) & x(620) & x(647) & x(648) & x(649) & x(652) & x(674) & x(676) & x(692) & x(693) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(732) & x(739) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(748);
    y(134) <= not(p134_out);
    p134 : perceptron
        Generic map (
            WEIGHTS => "0000000000000000000000000000000000000000000000000001111110010111111011011101000000000000000000000000000111111111111111111",
            SHIFT => 4,
            B => -648,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p134_in,
            y(0) => p134_out,
            y(1 to 17 - 1) => dummy134
        );


    p135_in <= x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(103) & x(104) & x(107) & x(108) & x(192) & x(199) & x(211) & x(220) & x(238) & x(239) & x(248) & x(249) & x(273) & x(274) & x(277) & x(299) & x(300) & x(305) & x(325) & x(326) & x(327) & x(342) & x(353) & x(354) & x(355) & x(360) & x(374) & x(380) & x(401) & x(402) & x(405) & x(407) & x(432) & x(433) & x(441) & x(460) & x(461) & x(463) & x(464) & x(473) & x(479) & x(487) & x(488) & x(489) & x(490) & x(491) & x(501) & x(502) & x(514) & x(516) & x(517) & x(518) & x(528) & x(529) & x(530) & x(556) & x(557) & x(558) & x(572) & x(573) & x(583) & x(584) & x(601) & x(610) & x(611) & x(612) & x(634) & x(637) & x(638) & x(639) & x(657) & x(660) & x(686) & x(688) & x(690) & x(695) & x(709) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(746) & x(747) & x(748);
    y(135) <= not(p135_out);
    p135 : perceptron
        Generic map (
            WEIGHTS => "00000000000000010010011111111111011100100111101111111111111111111111100110111111111111000000000000",
            SHIFT => 4,
            B => 20,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p135_in,
            y(0) => p135_out,
            y(1 to 16 - 1) => dummy135
        );


    p136_in <= x(77) & x(101) & x(102) & x(103) & x(104) & x(105) & x(106) & x(165) & x(193) & x(197) & x(198) & x(221) & x(226) & x(247) & x(248) & x(249) & x(275) & x(276) & x(277) & x(304) & x(309) & x(320) & x(330) & x(338) & x(347) & x(348) & x(349) & x(357) & x(362) & x(375) & x(376) & x(394) & x(397) & x(416) & x(444) & x(450) & x(473) & x(514) & x(515) & x(516) & x(535) & x(557) & x(647) & x(656) & x(657) & x(674) & x(675) & x(676) & x(677) & x(678) & x(716) & x(717) & x(718) & x(719) & x(721) & x(736) & x(737) & x(738) & x(739) & x(740) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(764) & x(766) & x(770) & x(771) & x(772) & x(773);
    y(136) <= not(p136_out);
    p136 : perceptron
        Generic map (
            WEIGHTS => "000000011101011111110100111011101111000010111111110000000000000000000000",
            SHIFT => 5,
            B => -288,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p136_in,
            y(0) => p136_out,
            y(1 to 17 - 1) => dummy136
        );


    p137_in <= x(37) & x(40) & x(41) & x(73) & x(74) & x(75) & x(77) & x(78) & x(79) & x(103) & x(104) & x(105) & x(106) & x(107) & x(133) & x(166) & x(193) & x(221) & x(247) & x(248) & x(249) & x(250) & x(275) & x(276) & x(277) & x(303) & x(306) & x(307) & x(334) & x(342) & x(358) & x(359) & x(361) & x(362) & x(367) & x(370) & x(371) & x(386) & x(387) & x(388) & x(390) & x(399) & x(414) & x(415) & x(416) & x(418) & x(433) & x(441) & x(442) & x(443) & x(446) & x(447) & x(473) & x(474) & x(500) & x(501) & x(502) & x(528) & x(529) & x(541) & x(556) & x(557) & x(558) & x(583) & x(584) & x(610) & x(611) & x(612) & x(638) & x(640);
    y(137) <= not(p137_out);
    p137 : perceptron
        Generic map (
            WEIGHTS => "1111111111111110000000000000011100011111011110011100000000000000000000",
            SHIFT => 5,
            B => -286,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p137_in,
            y(0) => p137_out,
            y(1 to 17 - 1) => dummy137
        );


    p138_in <= x(37) & x(39) & x(40) & x(41) & x(45) & x(46) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(73) & x(74) & x(75) & x(78) & x(79) & x(102) & x(103) & x(104) & x(105) & x(117) & x(118) & x(121) & x(165) & x(182) & x(193) & x(198) & x(207) & x(209) & x(214) & x(221) & x(234) & x(243) & x(244) & x(245) & x(247) & x(248) & x(249) & x(250) & x(275) & x(276) & x(277) & x(278) & x(294) & x(303) & x(304) & x(305) & x(306) & x(307) & x(333) & x(334) & x(347) & x(348) & x(358) & x(361) & x(362) & x(374) & x(376) & x(386) & x(387) & x(389) & x(390) & x(391) & x(400) & x(401) & x(402) & x(412) & x(414) & x(418) & x(427) & x(428) & x(429) & x(439) & x(440) & x(446) & x(450) & x(456) & x(457) & x(460) & x(474) & x(479) & x(488) & x(502) & x(507) & x(517) & x(534) & x(535) & x(545) & x(557) & x(563) & x(566) & x(574) & x(582) & x(591) & x(595) & x(597) & x(602) & x(619) & x(647) & x(655) & x(656) & x(657) & x(658) & x(675) & x(681) & x(682) & x(695) & x(719) & x(720) & x(721) & x(723) & x(747) & x(748) & x(749);
    y(138) <= not(p138_out);
    p138 : perceptron
        Generic map (
            WEIGHTS => "11111111111111111111110000001000000000000000010000000001001011000111110111110011000000100100010000100000000000000000",
            SHIFT => 4,
            B => -359,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p138_in,
            y(0) => p138_out,
            y(1 to 16 - 1) => dummy138
        );


    p139_in <= x(75) & x(78) & x(79) & x(104) & x(105) & x(106) & x(125) & x(126) & x(151) & x(152) & x(153) & x(154) & x(155) & x(166) & x(179) & x(180) & x(181) & x(182) & x(183) & x(184) & x(193) & x(194) & x(210) & x(211) & x(212) & x(220) & x(221) & x(222) & x(238) & x(248) & x(249) & x(250) & x(251) & x(276) & x(277) & x(278) & x(304) & x(305) & x(306) & x(309) & x(322) & x(333) & x(334) & x(337) & x(345) & x(349) & x(350) & x(351) & x(359) & x(360) & x(361) & x(362) & x(372) & x(373) & x(374) & x(377) & x(378) & x(387) & x(388) & x(390) & x(399) & x(400) & x(401) & x(402) & x(406) & x(414) & x(418) & x(425) & x(428) & x(429) & x(433) & x(446) & x(479) & x(507) & x(557) & x(566) & x(591) & x(624) & x(625) & x(652) & x(653) & x(694) & x(695) & x(704) & x(712) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(746) & x(747) & x(748) & x(749) & x(773);
    y(139) <= not(p139_out);
    p139 : perceptron
        Generic map (
            WEIGHTS => "00000011111111111111111111111111111111101110011100110001100100001010001111011111111011111111111110",
            SHIFT => 3,
            B => 310,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p139_in,
            y(0) => p139_out,
            y(1 to 15 - 1) => dummy139
        );


    p140_in <= x(35) & x(40) & x(63) & x(66) & x(67) & x(181) & x(182) & x(183) & x(184) & x(198) & x(210) & x(211) & x(212) & x(213) & x(239) & x(248) & x(249) & x(250) & x(276) & x(277) & x(278) & x(304) & x(306) & x(310) & x(311) & x(322) & x(334) & x(339) & x(344) & x(345) & x(346) & x(348) & x(349) & x(350) & x(361) & x(362) & x(371) & x(372) & x(373) & x(374) & x(375) & x(376) & x(377) & x(378) & x(450) & x(473) & x(502) & x(506) & x(507) & x(528) & x(530) & x(534) & x(535) & x(557) & x(558) & x(591) & x(619) & x(647) & x(648) & x(649) & x(674) & x(675) & x(676) & x(677) & x(693) & x(694) & x(695) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(732) & x(747) & x(748) & x(749) & x(769) & x(770) & x(773) & x(774);
    y(140) <= not(p140_out);
    p140 : perceptron
        Generic map (
            WEIGHTS => "0000000001000000000000011001111000001111100001100110011000000000000000000000001111",
            SHIFT => 4,
            B => -466,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p140_in,
            y(0) => p140_out,
            y(1 to 16 - 1) => dummy140
        );


    p141_in <= x(74) & x(75) & x(91) & x(104) & x(147) & x(175) & x(191) & x(192) & x(204) & x(210) & x(238) & x(242) & x(266) & x(267) & x(295) & x(320) & x(347) & x(348) & x(349) & x(374) & x(375) & x(390) & x(403) & x(404) & x(408) & x(418) & x(424) & x(431) & x(436) & x(439) & x(440) & x(443) & x(445) & x(446) & x(460) & x(463) & x(465) & x(473) & x(474) & x(479) & x(501) & x(502) & x(529) & x(548) & x(557) & x(576) & x(709) & x(710) & x(711) & x(712) & x(713) & x(714) & x(715) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(735) & x(736) & x(737) & x(738) & x(739) & x(740) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(748) & x(749);
    y(141) <= not(p141_out);
    p141 : perceptron
        Generic map (
            WEIGHTS => "0010000001111110000001000100000011000111111010111111111111111111111111111111",
            SHIFT => 4,
            B => 448,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p141_in,
            y(0) => p141_out,
            y(1 to 16 - 1) => dummy141
        );


    p142_in <= x(3) & x(25) & x(27) & x(34) & x(35) & x(36) & x(37) & x(38) & x(39) & x(40) & x(41) & x(43) & x(54) & x(58) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(79) & x(102) & x(103) & x(104) & x(105) & x(106) & x(107) & x(108) & x(118) & x(121) & x(151) & x(153) & x(168) & x(189) & x(192) & x(193) & x(194) & x(195) & x(215) & x(221) & x(222) & x(248) & x(249) & x(250) & x(268) & x(269) & x(276) & x(277) & x(278) & x(283) & x(295) & x(305) & x(306) & x(310) & x(311) & x(312) & x(317) & x(318) & x(319) & x(322) & x(323) & x(328) & x(329) & x(330) & x(331) & x(338) & x(339) & x(345) & x(349) & x(355) & x(357) & x(358) & x(359) & x(360) & x(362) & x(366) & x(379) & x(385) & x(386) & x(387) & x(388) & x(390) & x(392) & x(403) & x(405) & x(408) & x(414) & x(415) & x(418) & x(419) & x(431) & x(436) & x(446) & x(458) & x(473) & x(474) & x(479) & x(485) & x(486) & x(487) & x(500) & x(501) & x(502) & x(507) & x(513) & x(514) & x(515) & x(525) & x(528) & x(529) & x(530) & x(535) & x(536) & x(537) & x(543) & x(552) & x(555) & x(556) & x(557) & x(558) & x(563) & x(564) & x(566) & x(583) & x(584) & x(585) & x(591) & x(592) & x(597) & x(611) & x(612) & x(613) & x(615) & x(619) & x(620) & x(625) & x(638) & x(640) & x(648) & x(649) & x(650) & x(653) & x(677) & x(690) & x(691) & x(692) & x(693) & x(694) & x(695) & x(706) & x(707) & x(708) & x(709) & x(719) & x(720) & x(721) & x(722) & x(723) & x(727) & x(730) & x(748) & x(758) & x(759) & x(761) & x(764) & x(765) & x(766) & x(769) & x(770) & x(773) & x(774);
    y(142) <= not(p142_out);
    p142 : perceptron
        Generic map (
            WEIGHTS => "11111111111111111111111111111111111111100001000000000000000000000001110011110011111110011111011111101110100011100001110000000100000000000000000100000000001111110000111111111100000000",
            SHIFT => 4,
            B => -104,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p142_in,
            y(0) => p142_out,
            y(1 to 17 - 1) => dummy142
        );


    p143_in <= x(35) & x(37) & x(63) & x(66) & x(68) & x(92) & x(117) & x(132) & x(133) & x(145) & x(146) & x(152) & x(161) & x(171) & x(172) & x(173) & x(198) & x(226) & x(247) & x(248) & x(249) & x(254) & x(276) & x(277) & x(295) & x(305) & x(325) & x(326) & x(327) & x(330) & x(332) & x(333) & x(349) & x(350) & x(361) & x(366) & x(377) & x(378) & x(381) & x(382) & x(405) & x(406) & x(408) & x(409) & x(430) & x(433) & x(434) & x(436) & x(450) & x(451) & x(461) & x(464) & x(475) & x(478) & x(479) & x(506) & x(507) & x(517) & x(534) & x(535) & x(544) & x(562) & x(563) & x(583) & x(591) & x(611) & x(618) & x(619) & x(620) & x(647) & x(648) & x(704);
    y(143) <= not(p143_out);
    p143 : perceptron
        Generic map (
            WEIGHTS => "000000100111011100000000011111111110111111111111111111111011011010111110",
            SHIFT => 4,
            B => 167,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p143_in,
            y(0) => p143_out,
            y(1 to 16 - 1) => dummy143
        );


    p144_in <= x(2) & x(4) & x(6) & x(12) & x(25) & x(35) & x(36) & x(37) & x(38) & x(39) & x(40) & x(41) & x(42) & x(44) & x(55) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(79) & x(90) & x(91) & x(92) & x(93) & x(94) & x(95) & x(96) & x(97) & x(98) & x(99) & x(100) & x(101) & x(102) & x(103) & x(104) & x(105) & x(106) & x(110) & x(154) & x(183) & x(220) & x(221) & x(248) & x(249) & x(250) & x(269) & x(270) & x(276) & x(277) & x(297) & x(300) & x(305) & x(318) & x(322) & x(345) & x(350) & x(367) & x(370) & x(371) & x(378) & x(396) & x(397) & x(399) & x(406) & x(424) & x(425) & x(427) & x(445) & x(451) & x(456) & x(473) & x(479) & x(503) & x(507) & x(515) & x(524) & x(529) & x(534) & x(535) & x(542) & x(543) & x(544) & x(557) & x(563) & x(578) & x(591) & x(619) & x(647) & x(648) & x(652) & x(673) & x(674) & x(692) & x(693) & x(694) & x(719) & x(721) & x(722) & x(726) & x(759) & x(782);
    y(144) <= not(p144_out);
    p144 : perceptron
        Generic map (
            WEIGHTS => "000001111111110111111111111111111111111111111111110111111100110010101100100010001101101111111111111111101000000000",
            SHIFT => 4,
            B => 715,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p144_in,
            y(0) => p144_out,
            y(1 to 16 - 1) => dummy144
        );


    p145_in <= x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(91) & x(92) & x(104) & x(105) & x(106) & x(107) & x(108) & x(122) & x(123) & x(160) & x(161) & x(162) & x(171) & x(172) & x(173) & x(174) & x(176) & x(189) & x(190) & x(194) & x(199) & x(200) & x(201) & x(202) & x(220) & x(221) & x(222) & x(228) & x(248) & x(249) & x(250) & x(276) & x(277) & x(278) & x(297) & x(305) & x(306) & x(324) & x(325) & x(326) & x(327) & x(330) & x(332) & x(343) & x(360) & x(381) & x(398) & x(408) & x(409) & x(426) & x(436) & x(437) & x(438) & x(450) & x(464) & x(465) & x(478) & x(502) & x(506) & x(521) & x(528) & x(534) & x(535) & x(563) & x(568) & x(576) & x(583) & x(584) & x(591) & x(596) & x(597) & x(598) & x(611) & x(618) & x(619) & x(638) & x(640) & x(647) & x(648) & x(675) & x(676) & x(677) & x(679) & x(706) & x(714) & x(773);
    y(145) <= not(p145_out);
    p145 : perceptron
        Generic map (
            WEIGHTS => "11111111000000011100000111000011101111110110000001001001000000010010001011011110011000000000",
            SHIFT => 4,
            B => -96,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p145_in,
            y(0) => p145_out,
            y(1 to 16 - 1) => dummy145
        );


    p146_in <= x(44) & x(71) & x(72) & x(74) & x(75) & x(91) & x(93) & x(94) & x(102) & x(108) & x(136) & x(154) & x(155) & x(171) & x(199) & x(293) & x(305) & x(327) & x(342) & x(354) & x(371) & x(373) & x(374) & x(397) & x(405) & x(432) & x(433) & x(441) & x(442) & x(450) & x(473) & x(488) & x(490) & x(492) & x(501) & x(502) & x(506) & x(518) & x(528) & x(529) & x(530) & x(556) & x(557) & x(558) & x(571) & x(572) & x(573) & x(582) & x(583) & x(584) & x(602) & x(609) & x(610) & x(611) & x(612) & x(634) & x(635) & x(636) & x(637) & x(638) & x(639) & x(665) & x(675) & x(677) & x(679) & x(697) & x(706) & x(707) & x(708) & x(709) & x(712) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(746) & x(747) & x(748);
    y(146) <= not(p146_out);
    p146 : perceptron
        Generic map (
            WEIGHTS => "1000011100011000110100001110001111110111111100011101111111111100010000000000000000",
            SHIFT => 4,
            B => -165,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p146_in,
            y(0) => p146_out,
            y(1 to 16 - 1) => dummy146
        );


    p147_in <= x(0) & x(1) & x(2) & x(3) & x(4) & x(5) & x(6) & x(7) & x(8) & x(9) & x(10) & x(11) & x(12) & x(15) & x(16) & x(17) & x(18) & x(19) & x(20) & x(21) & x(22) & x(23) & x(24) & x(25) & x(26) & x(27) & x(28) & x(29) & x(30) & x(31) & x(32) & x(33) & x(40) & x(46) & x(52) & x(53) & x(54) & x(55) & x(56) & x(57) & x(58) & x(59) & x(61) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(79) & x(82) & x(83) & x(84) & x(85) & x(87) & x(88) & x(103) & x(104) & x(105) & x(106) & x(107) & x(108) & x(110) & x(111) & x(112) & x(113) & x(115) & x(125) & x(126) & x(127) & x(128) & x(129) & x(139) & x(140) & x(141) & x(142) & x(151) & x(153) & x(154) & x(155) & x(156) & x(167) & x(168) & x(169) & x(171) & x(172) & x(193) & x(196) & x(197) & x(199) & x(200) & x(220) & x(221) & x(248) & x(249) & x(262) & x(276) & x(277) & x(278) & x(304) & x(305) & x(306) & x(316) & x(319) & x(320) & x(321) & x(333) & x(334) & x(347) & x(348) & x(349) & x(353) & x(354) & x(361) & x(364) & x(375) & x(376) & x(377) & x(381) & x(392) & x(409) & x(419) & x(420) & x(436) & x(446) & x(448) & x(449) & x(450) & x(454) & x(464) & x(468) & x(473) & x(474) & x(476) & x(478) & x(481) & x(496) & x(501) & x(502) & x(503) & x(504) & x(506) & x(507) & x(518) & x(523) & x(524) & x(528) & x(529) & x(532) & x(534) & x(535) & x(542) & x(543) & x(544) & x(550) & x(551) & x(552) & x(556) & x(557) & x(558) & x(560) & x(563) & x(569) & x(570) & x(571) & x(572) & x(584) & x(587) & x(588) & x(598) & x(611) & x(612) & x(615) & x(616) & x(617) & x(638) & x(643) & x(644) & x(645) & x(647) & x(648) & x(671) & x(672) & x(673) & x(675) & x(676) & x(677) & x(679) & x(680) & x(681) & x(693) & x(698) & x(699) & x(700) & x(701) & x(702) & x(706) & x(707) & x(708) & x(709) & x(710) & x(714) & x(721) & x(725) & x(726) & x(727) & x(728) & x(729) & x(730) & x(731) & x(735) & x(736) & x(746) & x(749) & x(750) & x(752) & x(753) & x(754) & x(755) & x(756) & x(757) & x(758) & x(759) & x(760) & x(766) & x(767) & x(769) & x(770) & x(772) & x(773) & x(779) & x(780) & x(781) & x(782) & x(783);
    y(147) <= not(p147_out);
    p147 : perceptron
        Generic map (
            WEIGHTS => "111111111111111111111111111111110011111111100000000011111100000011111111111111111111110001000000000000000000000000001000010110111010111101111110011111100111111111101111111111111111100111000000011111000000011111110000011111111100000011111",
            SHIFT => 3,
            B => 637,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p147_in,
            y(0) => p147_out,
            y(1 to 17 - 1) => dummy147
        );


    p148_in <= x(35) & x(36) & x(37) & x(38) & x(39) & x(40) & x(41) & x(44) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(75) & x(76) & x(79) & x(90) & x(91) & x(92) & x(93) & x(94) & x(95) & x(96) & x(136) & x(145) & x(155) & x(171) & x(172) & x(173) & x(182) & x(197) & x(199) & x(200) & x(201) & x(228) & x(248) & x(249) & x(276) & x(291) & x(296) & x(297) & x(299) & x(301) & x(322) & x(323) & x(324) & x(325) & x(326) & x(327) & x(332) & x(333) & x(334) & x(350) & x(351) & x(361) & x(381) & x(402) & x(409) & x(422) & x(430) & x(436) & x(437) & x(450) & x(458) & x(473) & x(474) & x(478) & x(500) & x(501) & x(502) & x(506) & x(507) & x(511) & x(513) & x(514) & x(515) & x(523) & x(525) & x(526) & x(528) & x(529) & x(534) & x(535) & x(538) & x(539) & x(541) & x(542) & x(543) & x(544) & x(549) & x(557) & x(563) & x(568) & x(571) & x(582) & x(584) & x(595) & x(598) & x(608) & x(610) & x(611) & x(612) & x(618) & x(638) & x(640) & x(647) & x(648) & x(675) & x(676) & x(677) & x(679) & x(732) & x(736) & x(737);
    y(148) <= not(p148_out);
    p148 : perceptron
        Generic map (
            WEIGHTS => "0000000000000000000000000001101110111110000111111111111111110110111000100011000000000110000000010000000000100111111011",
            SHIFT => 4,
            B => -234,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p148_in,
            y(0) => p148_out,
            y(1 to 17 - 1) => dummy148
        );


    p149_in <= x(1) & x(3) & x(6) & x(7) & x(16) & x(18) & x(20) & x(21) & x(22) & x(23) & x(24) & x(27) & x(29) & x(30) & x(32) & x(41) & x(44) & x(52) & x(54) & x(55) & x(57) & x(58) & x(61) & x(74) & x(82) & x(88) & x(93) & x(94) & x(96) & x(108) & x(112) & x(115) & x(119) & x(121) & x(122) & x(141) & x(142) & x(164) & x(165) & x(166) & x(167) & x(168) & x(192) & x(193) & x(194) & x(195) & x(220) & x(221) & x(222) & x(248) & x(249) & x(250) & x(251) & x(276) & x(277) & x(278) & x(283) & x(292) & x(305) & x(306) & x(310) & x(311) & x(312) & x(328) & x(329) & x(330) & x(331) & x(333) & x(334) & x(338) & x(339) & x(340) & x(345) & x(357) & x(358) & x(359) & x(360) & x(362) & x(364) & x(366) & x(367) & x(385) & x(386) & x(387) & x(388) & x(390) & x(414) & x(416) & x(418) & x(419) & x(423) & x(445) & x(446) & x(447) & x(448) & x(451) & x(473) & x(474) & x(475) & x(479) & x(484) & x(487) & x(500) & x(501) & x(502) & x(507) & x(509) & x(510) & x(513) & x(515) & x(528) & x(529) & x(530) & x(531) & x(535) & x(537) & x(538) & x(555) & x(556) & x(557) & x(558) & x(563) & x(566) & x(567) & x(583) & x(584) & x(585) & x(587) & x(588) & x(591) & x(595) & x(596) & x(610) & x(611) & x(612) & x(613) & x(616) & x(619) & x(620) & x(625) & x(636) & x(638) & x(639) & x(640) & x(643) & x(644) & x(645) & x(671) & x(690) & x(691) & x(692) & x(693) & x(694) & x(695) & x(698) & x(700) & x(701) & x(702) & x(707) & x(708) & x(710) & x(711) & x(712) & x(719) & x(720) & x(721) & x(722) & x(725) & x(729) & x(730) & x(752) & x(753) & x(755) & x(757) & x(760) & x(761) & x(764) & x(765) & x(766) & x(767) & x(768) & x(769) & x(770) & x(771) & x(772) & x(773) & x(774) & x(780);
    y(149) <= not(p149_out);
    p149 : perceptron
        Generic map (
            WEIGHTS => "11111111111111110111111111000111000110001100000000000000010000011110000011111010011110110100001000001100000011000000000000000001100000001000000011111111111111000001111111111110000000000001",
            SHIFT => 4,
            B => -428,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p149_in,
            y(0) => p149_out,
            y(1 to 17 - 1) => dummy149
        );


    p150_in <= x(9) & x(17) & x(32) & x(34) & x(35) & x(37) & x(40) & x(41) & x(63) & x(64) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(79) & x(102) & x(103) & x(104) & x(105) & x(106) & x(107) & x(138) & x(139) & x(140) & x(165) & x(166) & x(192) & x(193) & x(194) & x(218) & x(219) & x(220) & x(221) & x(222) & x(231) & x(232) & x(234) & x(246) & x(247) & x(248) & x(249) & x(250) & x(257) & x(258) & x(259) & x(260) & x(264) & x(270) & x(271) & x(274) & x(275) & x(276) & x(277) & x(278) & x(283) & x(284) & x(304) & x(305) & x(306) & x(310) & x(311) & x(312) & x(320) & x(333) & x(334) & x(338) & x(339) & x(350) & x(357) & x(358) & x(359) & x(362) & x(366) & x(367) & x(383) & x(386) & x(387) & x(390) & x(391) & x(406) & x(414) & x(418) & x(429) & x(434) & x(446) & x(457) & x(458) & x(473) & x(474) & x(479) & x(484) & x(500) & x(501) & x(502) & x(515) & x(528) & x(529) & x(556) & x(557) & x(574) & x(584) & x(587) & x(644) & x(656) & x(657) & x(658) & x(659) & x(660) & x(671) & x(681) & x(691) & x(692) & x(693) & x(694) & x(695) & x(708) & x(719) & x(720) & x(721) & x(722) & x(727) & x(730) & x(743) & x(755) & x(761) & x(763) & x(764) & x(766) & x(769) & x(770) & x(771) & x(773) & x(774);
    y(150) <= not(p150_out);
    p150 : perceptron
        Generic map (
            WEIGHTS => "1111111111111111111111111111110110000000000000000000000000000000000000000000111100011100110110110001000100001011000001011111011111101000000000",
            SHIFT => 4,
            B => -240,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p150_in,
            y(0) => p150_out,
            y(1 to 17 - 1) => dummy150
        );


    p151_in <= x(34) & x(35) & x(36) & x(37) & x(38) & x(39) & x(40) & x(41) & x(43) & x(45) & x(46) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(79) & x(99) & x(100) & x(102) & x(103) & x(104) & x(105) & x(106) & x(107) & x(108) & x(133) & x(147) & x(161) & x(162) & x(174) & x(175) & x(182) & x(190) & x(210) & x(248) & x(269) & x(276) & x(297) & x(299) & x(301) & x(311) & x(320) & x(323) & x(324) & x(327) & x(328) & x(333) & x(338) & x(347) & x(348) & x(353) & x(354) & x(355) & x(359) & x(366) & x(381) & x(385) & x(386) & x(387) & x(388) & x(390) & x(401) & x(402) & x(406) & x(414) & x(415) & x(416) & x(418) & x(433) & x(435) & x(436) & x(441) & x(444) & x(446) & x(460) & x(463) & x(464) & x(468) & x(469) & x(473) & x(474) & x(475) & x(491) & x(495) & x(501) & x(502) & x(528) & x(529) & x(530) & x(542) & x(543) & x(544) & x(556) & x(557) & x(558) & x(584) & x(585) & x(601) & x(602) & x(612) & x(675) & x(721) & x(722) & x(723) & x(765) & x(770) & x(773);
    y(151) <= not(p151_out);
    p151 : perceptron
        Generic map (
            WEIGHTS => "111111111111111111111111111111111111111011000101010000100000011000100111101101110000110000110000100000111000001101111000",
            SHIFT => 4,
            B => 359,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p151_in,
            y(0) => p151_out,
            y(1 to 17 - 1) => dummy151
        );


    p152_in <= x(35) & x(36) & x(37) & x(38) & x(39) & x(40) & x(41) & x(44) & x(45) & x(46) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(79) & x(90) & x(91) & x(92) & x(93) & x(94) & x(99) & x(100) & x(101) & x(102) & x(103) & x(104) & x(105) & x(106) & x(131) & x(146) & x(171) & x(172) & x(198) & x(226) & x(244) & x(248) & x(249) & x(250) & x(254) & x(276) & x(277) & x(282) & x(298) & x(305) & x(309) & x(310) & x(314) & x(338) & x(339) & x(340) & x(360) & x(366) & x(367) & x(378) & x(394) & x(397) & x(400) & x(401) & x(403) & x(406) & x(417) & x(424) & x(425) & x(426) & x(427) & x(445) & x(446) & x(450) & x(453) & x(454) & x(466) & x(481) & x(515) & x(517) & x(534) & x(544) & x(592) & x(606) & x(620) & x(647) & x(648) & x(674) & x(675) & x(706) & x(707) & x(708) & x(709) & x(710) & x(711) & x(712) & x(713) & x(714) & x(715) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(735) & x(736) & x(737) & x(738) & x(739) & x(740) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(750) & x(764) & x(765) & x(766) & x(768) & x(769) & x(770) & x(771) & x(772) & x(773) & x(774);
    y(152) <= not(p152_out);
    p152 : perceptron
        Generic map (
            WEIGHTS => "00000000000000000000000000000000000000000011100100000001000000010000111100111101111110010111111100000000000000000000000000000000000000000",
            SHIFT => 4,
            B => -1684,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p152_in,
            y(0) => p152_out,
            y(1 to 17 - 1) => dummy152
        );


    p153_in <= x(198) & x(309) & x(322) & x(323) & x(338) & x(339) & x(347) & x(360) & x(366) & x(367) & x(375) & x(387) & x(388) & x(401) & x(403) & x(418) & x(425) & x(450) & x(472) & x(647) & x(675) & x(708) & x(712) & x(717) & x(718) & x(719) & x(720) & x(721) & x(735) & x(736) & x(737) & x(739) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(750) & x(764) & x(770) & x(773);
    y(153) <= not(p153_out);
    p153 : perceptron
        Generic map (
            WEIGHTS => "0000001100111110111110000000000000000000000",
            SHIFT => 5,
            B => -776,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p153_in,
            y(0) => p153_out,
            y(1 to 16 - 1) => dummy153
        );


    p154_in <= x(0) & x(1) & x(2) & x(3) & x(4) & x(5) & x(6) & x(7) & x(8) & x(9) & x(10) & x(11) & x(12) & x(15) & x(16) & x(17) & x(18) & x(19) & x(20) & x(21) & x(22) & x(23) & x(24) & x(25) & x(26) & x(27) & x(28) & x(29) & x(30) & x(31) & x(32) & x(33) & x(44) & x(52) & x(53) & x(54) & x(55) & x(56) & x(57) & x(58) & x(59) & x(61) & x(76) & x(82) & x(83) & x(84) & x(85) & x(87) & x(88) & x(93) & x(94) & x(96) & x(110) & x(111) & x(112) & x(113) & x(115) & x(139) & x(140) & x(141) & x(142) & x(165) & x(167) & x(168) & x(169) & x(193) & x(196) & x(197) & x(210) & x(219) & x(220) & x(221) & x(247) & x(248) & x(249) & x(250) & x(275) & x(276) & x(294) & x(295) & x(303) & x(304) & x(319) & x(320) & x(323) & x(330) & x(332) & x(334) & x(338) & x(342) & x(347) & x(348) & x(349) & x(361) & x(362) & x(364) & x(370) & x(376) & x(378) & x(390) & x(392) & x(419) & x(420) & x(445) & x(447) & x(448) & x(449) & x(473) & x(474) & x(476) & x(502) & x(503) & x(504) & x(514) & x(532) & x(541) & x(557) & x(560) & x(587) & x(588) & x(615) & x(616) & x(617) & x(643) & x(644) & x(645) & x(656) & x(657) & x(658) & x(671) & x(672) & x(673) & x(694) & x(698) & x(699) & x(700) & x(701) & x(702) & x(716) & x(718) & x(719) & x(720) & x(721) & x(722) & x(725) & x(726) & x(727) & x(728) & x(729) & x(730) & x(731) & x(739) & x(742) & x(746) & x(747) & x(748) & x(752) & x(753) & x(754) & x(755) & x(756) & x(757) & x(758) & x(759) & x(760) & x(773) & x(774) & x(779) & x(780) & x(781) & x(782) & x(783);
    y(154) <= not(p154_out);
    p154 : perceptron
        Generic map (
            WEIGHTS => "0000000000000000000000000000000010000000001000000111000000000100010101111111110011110111101111100101000110011010010110000000001110000000000000000000000000000000000001100000",
            SHIFT => 5,
            B => -1991,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p154_in,
            y(0) => p154_out,
            y(1 to 18 - 1) => dummy154
        );


    p155_in <= x(7) & x(8) & x(9) & x(24) & x(26) & x(39) & x(42) & x(43) & x(44) & x(52) & x(58) & x(59) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(76) & x(77) & x(78) & x(79) & x(84) & x(85) & x(90) & x(91) & x(92) & x(93) & x(94) & x(95) & x(96) & x(104) & x(105) & x(106) & x(111) & x(113) & x(142) & x(167) & x(168) & x(183) & x(193) & x(194) & x(220) & x(221) & x(248) & x(249) & x(250) & x(255) & x(256) & x(276) & x(277) & x(282) & x(283) & x(284) & x(297) & x(305) & x(306) & x(310) & x(333) & x(334) & x(348) & x(349) & x(362) & x(364) & x(376) & x(377) & x(390) & x(392) & x(420) & x(433) & x(445) & x(451) & x(454) & x(473) & x(479) & x(507) & x(511) & x(535) & x(545) & x(556) & x(563) & x(583) & x(588) & x(591) & x(612) & x(615) & x(619) & x(645) & x(652) & x(655) & x(656) & x(700) & x(708) & x(712) & x(713) & x(720) & x(721) & x(725) & x(735) & x(736) & x(737) & x(738) & x(739) & x(742) & x(753) & x(759) & x(760) & x(769) & x(771) & x(772) & x(779) & x(782);
    y(155) <= not(p155_out);
    p155 : perceptron
        Generic map (
            WEIGHTS => "000001111000111111111111111001111111111000001111111100110000110111110111001110111010010010010111000011000000000000000",
            SHIFT => 5,
            B => 212,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p155_in,
            y(0) => p155_out,
            y(1 to 17 - 1) => dummy155
        );


    p156_in <= x(3) & x(5) & x(9) & x(15) & x(17) & x(18) & x(21) & x(30) & x(33) & x(84) & x(87) & x(93) & x(94) & x(110) & x(138) & x(142) & x(164) & x(165) & x(166) & x(192) & x(193) & x(194) & x(217) & x(220) & x(221) & x(222) & x(247) & x(248) & x(249) & x(250) & x(251) & x(276) & x(277) & x(278) & x(295) & x(304) & x(305) & x(306) & x(333) & x(334) & x(340) & x(350) & x(358) & x(359) & x(360) & x(361) & x(362) & x(367) & x(376) & x(386) & x(387) & x(388) & x(390) & x(392) & x(397) & x(411) & x(412) & x(414) & x(415) & x(416) & x(418) & x(419) & x(425) & x(427) & x(433) & x(439) & x(445) & x(446) & x(451) & x(454) & x(456) & x(457) & x(460) & x(461) & x(473) & x(474) & x(476) & x(479) & x(501) & x(502) & x(507) & x(528) & x(529) & x(535) & x(556) & x(557) & x(563) & x(584) & x(591) & x(612) & x(616) & x(619) & x(640) & x(643) & x(647) & x(695) & x(704) & x(709) & x(710) & x(712) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(724) & x(741) & x(746) & x(747) & x(748) & x(749) & x(750) & x(759) & x(783);
    y(156) <= not(p156_out);
    p156 : perceptron
        Generic map (
            WEIGHTS => "11111111111001010000000000000000001000000011100001110111111101110100011100001000000000000010010010000000000000000011",
            SHIFT => 4,
            B => -736,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p156_in,
            y(0) => p156_out,
            y(1 to 17 - 1) => dummy156
        );


    p157_in <= x(2) & x(5) & x(7) & x(9) & x(20) & x(23) & x(26) & x(27) & x(28) & x(29) & x(30) & x(31) & x(32) & x(33) & x(40) & x(44) & x(52) & x(53) & x(55) & x(58) & x(63) & x(64) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(76) & x(77) & x(78) & x(79) & x(82) & x(84) & x(88) & x(91) & x(93) & x(94) & x(95) & x(96) & x(97) & x(98) & x(99) & x(100) & x(101) & x(102) & x(103) & x(104) & x(105) & x(106) & x(110) & x(111) & x(112) & x(115) & x(122) & x(139) & x(146) & x(147) & x(151) & x(153) & x(154) & x(167) & x(169) & x(196) & x(198) & x(226) & x(289) & x(290) & x(305) & x(314) & x(315) & x(342) & x(343) & x(344) & x(345) & x(353) & x(361) & x(362) & x(364) & x(392) & x(445) & x(448) & x(450) & x(468) & x(470) & x(472) & x(473) & x(479) & x(497) & x(501) & x(502) & x(507) & x(522) & x(526) & x(528) & x(529) & x(534) & x(535) & x(550) & x(551) & x(553) & x(556) & x(557) & x(558) & x(563) & x(564) & x(578) & x(584) & x(591) & x(592) & x(602) & x(612) & x(616) & x(618) & x(619) & x(620) & x(644) & x(647) & x(648) & x(657) & x(660) & x(671) & x(674) & x(675) & x(676) & x(677) & x(691) & x(692) & x(698) & x(699) & x(701) & x(702) & x(725) & x(727) & x(728) & x(729) & x(732) & x(756) & x(757) & x(779) & x(780) & x(783);
    y(157) <= not(p157_out);
    p157 : perceptron
        Generic map (
            WEIGHTS => "1111111111111100111100000000000000011100000000000000011110100000111111101111111111101000000000000000000000000000000100010011100001111111111011111",
            SHIFT => 4,
            B => -238,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p157_in,
            y(0) => p157_out,
            y(1 to 17 - 1) => dummy157
        );


    p158_in <= x(45) & x(108) & x(135) & x(163) & x(164) & x(165) & x(182) & x(183) & x(184) & x(191) & x(192) & x(193) & x(194) & x(195) & x(197) & x(210) & x(211) & x(212) & x(219) & x(220) & x(221) & x(222) & x(237) & x(238) & x(239) & x(240) & x(247) & x(248) & x(249) & x(250) & x(276) & x(277) & x(278) & x(301) & x(302) & x(303) & x(304) & x(305) & x(326) & x(327) & x(328) & x(329) & x(330) & x(331) & x(332) & x(347) & x(356) & x(357) & x(358) & x(359) & x(360) & x(390) & x(400) & x(418) & x(450) & x(487) & x(501) & x(507) & x(513) & x(514) & x(515) & x(535) & x(542) & x(543) & x(563) & x(648) & x(675) & x(676) & x(677) & x(692) & x(693) & x(695) & x(703) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(740) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(748) & x(749);
    y(158) <= not(p158_out);
    p158 : perceptron
        Generic map (
            WEIGHTS => "1011110001111110001111000011111110000100000001000000101001000100111110001000000000000000000",
            SHIFT => 4,
            B => -94,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p158_in,
            y(0) => p158_out,
            y(1 to 16 - 1) => dummy158
        );


    p159_in <= x(35) & x(36) & x(37) & x(38) & x(39) & x(40) & x(41) & x(45) & x(46) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(79) & x(101) & x(102) & x(103) & x(104) & x(105) & x(106) & x(107) & x(108) & x(125) & x(126) & x(127) & x(182) & x(183) & x(184) & x(192) & x(193) & x(200) & x(210) & x(211) & x(248) & x(249) & x(250) & x(277) & x(304) & x(330) & x(331) & x(332) & x(338) & x(354) & x(355) & x(358) & x(359) & x(360) & x(366) & x(368) & x(371) & x(374) & x(378) & x(386) & x(387) & x(388) & x(398) & x(399) & x(400) & x(402) & x(405) & x(406) & x(413) & x(414) & x(415) & x(418) & x(426) & x(427) & x(433) & x(439) & x(440) & x(441) & x(446) & x(450) & x(460) & x(461) & x(467) & x(468) & x(487) & x(488) & x(501) & x(502) & x(528) & x(529) & x(530) & x(556) & x(557) & x(584) & x(665) & x(666) & x(676) & x(693) & x(694);
    y(159) <= not(p159_out);
    p159 : perceptron
        Generic map (
            WEIGHTS => "000000000000000000000000000000000001111111101111110000011000010010000000110001001000101100111111111111011",
            SHIFT => 4,
            B => -414,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p159_in,
            y(0) => p159_out,
            y(1 to 16 - 1) => dummy159
        );


    p160_in <= x(0) & x(1) & x(2) & x(3) & x(4) & x(5) & x(6) & x(7) & x(8) & x(9) & x(10) & x(11) & x(12) & x(15) & x(16) & x(17) & x(18) & x(19) & x(20) & x(21) & x(22) & x(23) & x(24) & x(25) & x(26) & x(27) & x(28) & x(29) & x(30) & x(31) & x(32) & x(33) & x(52) & x(53) & x(54) & x(55) & x(56) & x(57) & x(58) & x(59) & x(61) & x(67) & x(69) & x(70) & x(82) & x(83) & x(84) & x(85) & x(87) & x(88) & x(91) & x(93) & x(94) & x(97) & x(98) & x(110) & x(111) & x(112) & x(113) & x(115) & x(139) & x(140) & x(141) & x(142) & x(167) & x(168) & x(169) & x(182) & x(183) & x(190) & x(196) & x(197) & x(210) & x(211) & x(249) & x(250) & x(276) & x(277) & x(278) & x(305) & x(306) & x(333) & x(334) & x(350) & x(351) & x(360) & x(364) & x(377) & x(378) & x(388) & x(390) & x(392) & x(398) & x(400) & x(406) & x(414) & x(416) & x(418) & x(419) & x(420) & x(426) & x(445) & x(446) & x(448) & x(449) & x(473) & x(474) & x(475) & x(476) & x(479) & x(487) & x(501) & x(502) & x(503) & x(504) & x(515) & x(529) & x(532) & x(557) & x(560) & x(587) & x(588) & x(615) & x(616) & x(617) & x(643) & x(644) & x(645) & x(671) & x(672) & x(673) & x(675) & x(698) & x(699) & x(700) & x(701) & x(702) & x(709) & x(711) & x(712) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(725) & x(726) & x(727) & x(728) & x(729) & x(730) & x(731) & x(740) & x(741) & x(742) & x(744) & x(745) & x(746) & x(747) & x(748) & x(749) & x(752) & x(753) & x(754) & x(755) & x(756) & x(757) & x(758) & x(759) & x(760) & x(779) & x(780) & x(781) & x(782) & x(783);
    y(160) <= not(p160_out);
    p160 : perceptron
        Generic map (
            WEIGHTS => "0000000000000000000000000000000000000000011100000011111000000000000110001111111111111001101000100100011001110111100110100000000000000000011111111111000000011111111100000000000000",
            SHIFT => 5,
            B => -499,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p160_in,
            y(0) => p160_out,
            y(1 to 18 - 1) => dummy160
        );


    p161_in <= x(71) & x(72) & x(73) & x(74) & x(103) & x(104) & x(105) & x(106) & x(127) & x(129) & x(135) & x(136) & x(163) & x(164) & x(165) & x(166) & x(189) & x(191) & x(192) & x(193) & x(194) & x(199) & x(201) & x(207) & x(220) & x(221) & x(222) & x(245) & x(247) & x(248) & x(249) & x(250) & x(266) & x(276) & x(277) & x(278) & x(293) & x(294) & x(305) & x(320) & x(321) & x(329) & x(331) & x(333) & x(334) & x(340) & x(342) & x(347) & x(348) & x(349) & x(376) & x(377) & x(380) & x(381) & x(409) & x(416) & x(422) & x(423) & x(450) & x(454) & x(481) & x(501) & x(502) & x(507) & x(514) & x(518) & x(529) & x(535) & x(543) & x(545) & x(546) & x(557) & x(563) & x(584) & x(585) & x(611) & x(612) & x(618) & x(655) & x(656) & x(675) & x(676) & x(677) & x(678) & x(679);
    y(161) <= not(p161_out);
    p161 : perceptron
        Generic map (
            WEIGHTS => "0000000011000000000000000000000010001100011000000000000000011110111011110111100000000",
            SHIFT => 4,
            B => -679,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p161_in,
            y(0) => p161_out,
            y(1 to 16 - 1) => dummy161
        );


    p162_in <= x(64) & x(94) & x(118) & x(146) & x(152) & x(153) & x(154) & x(155) & x(156) & x(157) & x(173) & x(192) & x(200) & x(249) & x(256) & x(267) & x(277) & x(295) & x(301) & x(302) & x(303) & x(304) & x(311) & x(317) & x(329) & x(330) & x(331) & x(332) & x(333) & x(338) & x(342) & x(346) & x(361) & x(362) & x(369) & x(370) & x(371) & x(372) & x(374) & x(389) & x(390) & x(396) & x(397) & x(399) & x(401) & x(406) & x(418) & x(433) & x(434) & x(437) & x(445) & x(446) & x(473) & x(474) & x(479) & x(501) & x(502) & x(507) & x(514) & x(529) & x(534) & x(535) & x(541) & x(554) & x(557) & x(558) & x(563) & x(580) & x(591) & x(607) & x(609) & x(619) & x(624) & x(647) & x(692) & x(693) & x(694) & x(718) & x(719) & x(720) & x(721) & x(722) & x(748);
    y(162) <= not(p162_out);
    p162 : perceptron
        Generic map (
            WEIGHTS => "10000000000101001000000100000011001111100111100001000000000000000000000000111111111",
            SHIFT => 4,
            B => -414,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p162_in,
            y(0) => p162_out,
            y(1 to 16 - 1) => dummy162
        );


    p163_in <= x(2) & x(9) & x(22) & x(44) & x(54) & x(57) & x(67) & x(91) & x(92) & x(93) & x(94) & x(95) & x(115) & x(121) & x(138) & x(165) & x(166) & x(192) & x(193) & x(194) & x(220) & x(221) & x(222) & x(248) & x(249) & x(250) & x(276) & x(277) & x(278) & x(300) & x(302) & x(305) & x(306) & x(329) & x(330) & x(331) & x(332) & x(333) & x(334) & x(357) & x(358) & x(359) & x(360) & x(362) & x(367) & x(370) & x(371) & x(378) & x(386) & x(387) & x(388) & x(390) & x(397) & x(414) & x(415) & x(416) & x(418) & x(424) & x(425) & x(427) & x(443) & x(444) & x(445) & x(446) & x(448) & x(451) & x(453) & x(454) & x(455) & x(461) & x(473) & x(474) & x(479) & x(484) & x(485) & x(501) & x(502) & x(507) & x(528) & x(529) & x(530) & x(535) & x(556) & x(557) & x(563) & x(584) & x(591) & x(619) & x(636) & x(700) & x(709) & x(710) & x(711) & x(712) & x(719) & x(720) & x(721) & x(722) & x(723) & x(726) & x(730) & x(737) & x(747) & x(748) & x(749) & x(759) & x(782);
    y(163) <= not(p163_out);
    p163 : perceptron
        Generic map (
            WEIGHTS => "11101100000010000000000000000110011110011110011011101111011111001011100001100000000000000100000000011000011",
            SHIFT => 4,
            B => -489,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p163_in,
            y(0) => p163_out,
            y(1 to 16 - 1) => dummy163
        );


    p164_in <= x(91) & x(92) & x(93) & x(171) & x(172) & x(197) & x(198) & x(200) & x(201) & x(213) & x(266) & x(272) & x(293) & x(294) & x(322) & x(347) & x(348) & x(350) & x(360) & x(375) & x(376) & x(380) & x(388) & x(397) & x(398) & x(399) & x(400) & x(414) & x(415) & x(416) & x(418) & x(425) & x(426) & x(427) & x(428) & x(429) & x(430) & x(431) & x(436) & x(443) & x(444) & x(450) & x(456) & x(466) & x(473) & x(474) & x(489) & x(501) & x(502) & x(506) & x(516) & x(517) & x(528) & x(529) & x(534) & x(535) & x(545) & x(557) & x(562) & x(563) & x(583) & x(584) & x(605) & x(611) & x(618) & x(638) & x(646) & x(647) & x(648) & x(674) & x(675) & x(676) & x(677) & x(678) & x(679) & x(713) & x(716) & x(718) & x(739) & x(741) & x(742) & x(744) & x(745) & x(746);
    y(164) <= not(p164_out);
    p164 : perceptron
        Generic map (
            WEIGHTS => "111000100010111001000000000000100000000000001111101111001100110101000000000111111111",
            SHIFT => 4,
            B => -140,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p164_in,
            y(0) => p164_out,
            y(1 to 16 - 1) => dummy164
        );


    p165_in <= x(2) & x(5) & x(6) & x(7) & x(8) & x(12) & x(16) & x(18) & x(20) & x(21) & x(23) & x(25) & x(29) & x(33) & x(35) & x(36) & x(37) & x(38) & x(39) & x(40) & x(41) & x(42) & x(44) & x(45) & x(46) & x(53) & x(54) & x(56) & x(57) & x(61) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(79) & x(85) & x(90) & x(91) & x(92) & x(93) & x(94) & x(95) & x(96) & x(97) & x(98) & x(99) & x(100) & x(101) & x(102) & x(103) & x(104) & x(105) & x(106) & x(107) & x(108) & x(110) & x(111) & x(136) & x(141) & x(152) & x(155) & x(163) & x(164) & x(165) & x(166) & x(167) & x(169) & x(182) & x(190) & x(192) & x(193) & x(196) & x(219) & x(220) & x(244) & x(247) & x(248) & x(249) & x(263) & x(276) & x(288) & x(290) & x(294) & x(307) & x(314) & x(317) & x(318) & x(319) & x(322) & x(323) & x(334) & x(344) & x(347) & x(349) & x(353) & x(366) & x(378) & x(420) & x(449) & x(450) & x(479) & x(496) & x(499) & x(507) & x(529) & x(535) & x(543) & x(544) & x(551) & x(557) & x(563) & x(564) & x(584) & x(587) & x(591) & x(592) & x(602) & x(612) & x(615) & x(619) & x(620) & x(643) & x(647) & x(648) & x(649) & x(657) & x(661) & x(671) & x(672) & x(674) & x(675) & x(676) & x(677) & x(678) & x(690) & x(691) & x(692) & x(693) & x(695) & x(699) & x(719) & x(721) & x(722) & x(727) & x(728) & x(729) & x(754) & x(756) & x(757) & x(758) & x(759) & x(760) & x(781);
    y(165) <= not(p165_out);
    p165 : perceptron
        Generic map (
            WEIGHTS => "0000000000000011111111111000001111111111111111110111111111111111111100001100000010000000000000010000011000001100111111111111110111101101110000111110000000000000000000",
            SHIFT => 4,
            B => 18,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p165_in,
            y(0) => p165_out,
            y(1 to 17 - 1) => dummy165
        );


    p166_in <= x(64) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(91) & x(93) & x(94) & x(102) & x(103) & x(104) & x(105) & x(106) & x(107) & x(108) & x(171) & x(172) & x(193) & x(197) & x(199) & x(200) & x(201) & x(219) & x(221) & x(227) & x(228) & x(247) & x(248) & x(249) & x(267) & x(275) & x(276) & x(277) & x(291) & x(294) & x(295) & x(296) & x(322) & x(323) & x(324) & x(405) & x(414) & x(415) & x(416) & x(432) & x(433) & x(441) & x(443) & x(446) & x(450) & x(460) & x(461) & x(473) & x(474) & x(487) & x(488) & x(489) & x(500) & x(501) & x(502) & x(506) & x(507) & x(514) & x(515) & x(516) & x(517) & x(518) & x(528) & x(529) & x(530) & x(534) & x(535) & x(542) & x(543) & x(556) & x(557) & x(558) & x(563) & x(583) & x(584) & x(610) & x(611) & x(612) & x(618) & x(637) & x(638) & x(639) & x(640) & x(647) & x(648) & x(649) & x(665) & x(667) & x(675) & x(676) & x(677) & x(678) & x(679) & x(697) & x(705) & x(706) & x(707) & x(708) & x(709) & x(718) & x(719) & x(720) & x(721) & x(735) & x(736) & x(737) & x(739) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(764) & x(765) & x(766) & x(770) & x(773);
    y(166) <= not(p166_out);
    p166 : perceptron
        Generic map (
            WEIGHTS => "011111111100011111111101111001100010000111111011100110100000000001100000000110000010000010000111001111101111111111111111111111111",
            SHIFT => 4,
            B => 407,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p166_in,
            y(0) => p166_out,
            y(1 to 17 - 1) => dummy166
        );


    p167_in <= x(35) & x(62) & x(68) & x(70) & x(78) & x(79) & x(96) & x(97) & x(99) & x(100) & x(101) & x(102) & x(105) & x(106) & x(108) & x(164) & x(165) & x(166) & x(191) & x(192) & x(193) & x(200) & x(219) & x(220) & x(221) & x(247) & x(248) & x(249) & x(250) & x(276) & x(277) & x(300) & x(305) & x(306) & x(309) & x(310) & x(326) & x(329) & x(333) & x(334) & x(338) & x(348) & x(349) & x(350) & x(358) & x(359) & x(366) & x(376) & x(377) & x(378) & x(405) & x(406) & x(432) & x(433) & x(434) & x(460) & x(461) & x(462) & x(529) & x(557) & x(638) & x(706) & x(707) & x(708) & x(709) & x(715) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(736) & x(737) & x(738) & x(739) & x(740) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(764) & x(766) & x(769) & x(770) & x(773) & x(774);
    y(167) <= not(p167_out);
    p167 : perceptron
        Generic map (
            WEIGHTS => "000000000000000111111011111111101100001101110001111111111100000000000000000000000000000000",
            SHIFT => 4,
            B => -507,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p167_in,
            y(0) => p167_out,
            y(1 to 16 - 1) => dummy167
        );


    p168_in <= x(1) & x(2) & x(5) & x(6) & x(7) & x(10) & x(11) & x(15) & x(17) & x(18) & x(20) & x(21) & x(22) & x(24) & x(26) & x(28) & x(33) & x(53) & x(54) & x(55) & x(57) & x(78) & x(79) & x(83) & x(84) & x(85) & x(88) & x(96) & x(101) & x(105) & x(106) & x(107) & x(108) & x(110) & x(112) & x(115) & x(118) & x(133) & x(135) & x(139) & x(151) & x(152) & x(153) & x(154) & x(155) & x(156) & x(162) & x(163) & x(164) & x(167) & x(168) & x(169) & x(171) & x(172) & x(173) & x(174) & x(175) & x(177) & x(178) & x(179) & x(180) & x(183) & x(184) & x(185) & x(192) & x(196) & x(197) & x(200) & x(209) & x(249) & x(254) & x(277) & x(297) & x(299) & x(300) & x(301) & x(302) & x(303) & x(304) & x(315) & x(317) & x(329) & x(330) & x(331) & x(332) & x(342) & x(343) & x(355) & x(358) & x(359) & x(360) & x(361) & x(370) & x(371) & x(376) & x(383) & x(384) & x(388) & x(389) & x(390) & x(399) & x(419) & x(420) & x(448) & x(450) & x(474) & x(476) & x(478) & x(479) & x(501) & x(502) & x(507) & x(514) & x(529) & x(534) & x(535) & x(540) & x(541) & x(545) & x(546) & x(551) & x(552) & x(553) & x(557) & x(562) & x(563) & x(565) & x(566) & x(567) & x(568) & x(569) & x(573) & x(584) & x(588) & x(590) & x(591) & x(593) & x(594) & x(595) & x(596) & x(615) & x(616) & x(618) & x(619) & x(620) & x(622) & x(623) & x(625) & x(626) & x(644) & x(647) & x(648) & x(654) & x(655) & x(656) & x(672) & x(673) & x(675) & x(717) & x(718) & x(719) & x(720) & x(721) & x(723) & x(725) & x(726) & x(745) & x(747) & x(748) & x(749) & x(753) & x(754) & x(758) & x(759) & x(781) & x(782);
    y(168) <= not(p168_out);
    p168 : perceptron
        Generic map (
            WEIGHTS => "11111111111111111111100111100000011101110000001111110000000000001100011100000001100001110000110110001111001000000000001100000000000101000000110000000100000110000000110000111111",
            SHIFT => 3,
            B => -116,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p168_in,
            y(0) => p168_out,
            y(1 to 16 - 1) => dummy168
        );


    p169_in <= x(34) & x(35) & x(37) & x(39) & x(40) & x(43) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(92) & x(118) & x(123) & x(125) & x(154) & x(164) & x(165) & x(166) & x(171) & x(172) & x(173) & x(174) & x(176) & x(178) & x(179) & x(184) & x(191) & x(192) & x(193) & x(194) & x(197) & x(199) & x(200) & x(201) & x(209) & x(220) & x(221) & x(222) & x(228) & x(248) & x(249) & x(250) & x(256) & x(276) & x(277) & x(278) & x(290) & x(291) & x(295) & x(296) & x(297) & x(298) & x(299) & x(300) & x(301) & x(302) & x(303) & x(305) & x(306) & x(310) & x(311) & x(315) & x(316) & x(317) & x(327) & x(329) & x(330) & x(331) & x(332) & x(334) & x(338) & x(342) & x(343) & x(344) & x(350) & x(359) & x(360) & x(378) & x(405) & x(422) & x(425) & x(446) & x(450) & x(453) & x(462) & x(474) & x(490) & x(501) & x(502) & x(529) & x(534) & x(535) & x(549) & x(550) & x(552) & x(556) & x(557) & x(558) & x(563) & x(581) & x(584) & x(591) & x(594) & x(595) & x(612) & x(619) & x(621) & x(622) & x(625) & x(647) & x(675) & x(676) & x(691) & x(692) & x(693) & x(694) & x(695) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(748) & x(749) & x(769);
    y(169) <= not(p169_out);
    p169 : perceptron
        Generic map (
            WEIGHTS => "11111111111111110000111000000001111000001110111011111000000000110011100000101111001100000101000000000000000000000000011111111111110",
            SHIFT => 4,
            B => -33,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p169_in,
            y(0) => p169_out,
            y(1 to 17 - 1) => dummy169
        );


    p170_in <= x(67) & x(68) & x(70) & x(77) & x(78) & x(79) & x(93) & x(94) & x(95) & x(96) & x(97) & x(101) & x(102) & x(103) & x(104) & x(105) & x(106) & x(107) & x(108) & x(121) & x(122) & x(192) & x(198) & x(221) & x(222) & x(248) & x(249) & x(263) & x(264) & x(276) & x(277) & x(292) & x(305) & x(309) & x(310) & x(322) & x(323) & x(329) & x(330) & x(333) & x(334) & x(338) & x(339) & x(349) & x(350) & x(351) & x(357) & x(366) & x(377) & x(378) & x(394) & x(406) & x(416) & x(424) & x(443) & x(445) & x(450) & x(473) & x(474) & x(487) & x(501) & x(502) & x(506) & x(514) & x(515) & x(528) & x(529) & x(530) & x(535) & x(556) & x(557) & x(584) & x(674) & x(675) & x(678) & x(707) & x(708) & x(709) & x(710) & x(711) & x(712) & x(714) & x(715) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(736) & x(737) & x(738) & x(739) & x(740) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(748) & x(750) & x(764) & x(765) & x(769) & x(770) & x(773) & x(774) & x(775);
    y(170) <= not(p170_out);
    p170 : perceptron
        Generic map (
            WEIGHTS => "00000000000000000000010111100110100110011001110011011110100000100000100011100000000000000000000000000000000000",
            SHIFT => 4,
            B => -953,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p170_in,
            y(0) => p170_out,
            y(1 to 16 - 1) => dummy170
        );


    p171_in <= x(36) & x(37) & x(45) & x(62) & x(63) & x(64) & x(65) & x(66) & x(68) & x(90) & x(91) & x(92) & x(93) & x(94) & x(107) & x(108) & x(164) & x(165) & x(172) & x(190) & x(191) & x(192) & x(193) & x(194) & x(199) & x(200) & x(218) & x(219) & x(220) & x(221) & x(222) & x(246) & x(247) & x(248) & x(249) & x(250) & x(267) & x(275) & x(276) & x(277) & x(291) & x(292) & x(294) & x(295) & x(296) & x(297) & x(298) & x(299) & x(301) & x(302) & x(309) & x(319) & x(320) & x(322) & x(323) & x(324) & x(325) & x(326) & x(327) & x(328) & x(329) & x(330) & x(331) & x(332) & x(338) & x(347) & x(348) & x(350) & x(351) & x(390) & x(446) & x(474) & x(475) & x(479) & x(507) & x(534) & x(535) & x(562) & x(563) & x(591) & x(619) & x(620) & x(646) & x(647) & x(648) & x(677) & x(720) & x(721) & x(739) & x(740) & x(741) & x(742) & x(743) & x(746) & x(747);
    y(171) <= not(p171_out);
    p171 : perceptron
        Generic map (
            WEIGHTS => "11111111111111001101111100111111111101111100000000011000000000000110000000000000000000000000000",
            SHIFT => 4,
            B => -103,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p171_in,
            y(0) => p171_out,
            y(1 to 16 - 1) => dummy171
        );


    p172_in <= x(0) & x(1) & x(2) & x(3) & x(4) & x(5) & x(6) & x(7) & x(8) & x(9) & x(10) & x(11) & x(12) & x(15) & x(16) & x(17) & x(18) & x(19) & x(20) & x(21) & x(22) & x(23) & x(24) & x(25) & x(26) & x(27) & x(28) & x(29) & x(30) & x(31) & x(32) & x(33) & x(37) & x(39) & x(40) & x(41) & x(46) & x(52) & x(53) & x(54) & x(55) & x(56) & x(57) & x(58) & x(59) & x(61) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(78) & x(79) & x(82) & x(83) & x(84) & x(85) & x(87) & x(88) & x(101) & x(102) & x(103) & x(104) & x(105) & x(110) & x(111) & x(112) & x(113) & x(115) & x(121) & x(139) & x(140) & x(141) & x(142) & x(146) & x(147) & x(165) & x(167) & x(168) & x(169) & x(175) & x(183) & x(186) & x(193) & x(196) & x(198) & x(199) & x(212) & x(226) & x(227) & x(237) & x(240) & x(247) & x(248) & x(249) & x(250) & x(262) & x(264) & x(271) & x(275) & x(276) & x(277) & x(278) & x(287) & x(288) & x(289) & x(290) & x(291) & x(302) & x(303) & x(307) & x(309) & x(310) & x(320) & x(322) & x(330) & x(331) & x(338) & x(339) & x(350) & x(361) & x(362) & x(364) & x(366) & x(367) & x(378) & x(386) & x(387) & x(389) & x(390) & x(392) & x(394) & x(401) & x(406) & x(414) & x(418) & x(419) & x(420) & x(434) & x(438) & x(446) & x(448) & x(449) & x(462) & x(468) & x(474) & x(476) & x(490) & x(500) & x(502) & x(503) & x(504) & x(510) & x(517) & x(532) & x(539) & x(540) & x(557) & x(560) & x(587) & x(588) & x(602) & x(603) & x(615) & x(616) & x(617) & x(643) & x(644) & x(645) & x(648) & x(656) & x(657) & x(658) & x(671) & x(672) & x(673) & x(698) & x(699) & x(700) & x(701) & x(702) & x(707) & x(709) & x(710) & x(711) & x(712) & x(713) & x(715) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(725) & x(726) & x(727) & x(728) & x(729) & x(730) & x(731) & x(736) & x(737) & x(738) & x(739) & x(740) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(748) & x(750) & x(752) & x(753) & x(754) & x(755) & x(756) & x(757) & x(758) & x(759) & x(760) & x(761) & x(764) & x(765) & x(766) & x(769) & x(770) & x(771) & x(773) & x(774) & x(779) & x(780) & x(781) & x(782) & x(783);
    y(172) <= not(p172_out);
    p172 : perceptron
        Generic map (
            WEIGHTS => "11111111111111111111111111111111111111111111111111111111111111111111111111111110111111011110001000000000000000000000000000001000010010011100101110111101111011001101100011111111111100011111111000000000000011111110000000000000011111111100000000011111",
            SHIFT => 4,
            B => -103,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p172_in,
            y(0) => p172_out,
            y(1 to 18 - 1) => dummy172
        );


    p173_in <= x(35) & x(38) & x(39) & x(40) & x(41) & x(43) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(78) & x(79) & x(89) & x(97) & x(98) & x(99) & x(105) & x(106) & x(107) & x(108) & x(162) & x(163) & x(164) & x(181) & x(182) & x(184) & x(190) & x(191) & x(192) & x(204) & x(209) & x(210) & x(211) & x(212) & x(218) & x(219) & x(220) & x(229) & x(231) & x(232) & x(237) & x(238) & x(239) & x(247) & x(248) & x(249) & x(250) & x(257) & x(266) & x(267) & x(277) & x(305) & x(328) & x(330) & x(331) & x(332) & x(333) & x(334) & x(347) & x(350) & x(412) & x(439) & x(440) & x(446) & x(462) & x(490) & x(502) & x(515) & x(517) & x(528) & x(530) & x(556) & x(584) & x(692) & x(693) & x(694) & x(695) & x(703) & x(712) & x(713) & x(714) & x(715) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(739) & x(740) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(748) & x(749);
    y(173) <= not(p173_out);
    p173 : perceptron
        Generic map (
            WEIGHTS => "11111111111111111111111111000111000011110000001110000011001111000100000001000001111011111111111111111111111",
            SHIFT => 4,
            B => 456,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p173_in,
            y(0) => p173_out,
            y(1 to 16 - 1) => dummy173
        );


    p174_in <= x(34) & x(35) & x(36) & x(37) & x(38) & x(39) & x(40) & x(41) & x(43) & x(45) & x(46) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(79) & x(102) & x(103) & x(104) & x(105) & x(106) & x(118) & x(192) & x(198) & x(199) & x(216) & x(226) & x(227) & x(248) & x(254) & x(255) & x(256) & x(266) & x(267) & x(268) & x(269) & x(270) & x(282) & x(283) & x(284) & x(294) & x(295) & x(296) & x(297) & x(309) & x(310) & x(311) & x(312) & x(326) & x(338) & x(339) & x(346) & x(347) & x(348) & x(349) & x(350) & x(352) & x(353) & x(354) & x(355) & x(359) & x(361) & x(362) & x(366) & x(370) & x(371) & x(374) & x(375) & x(376) & x(377) & x(378) & x(380) & x(381) & x(382) & x(386) & x(387) & x(390) & x(394) & x(405) & x(414) & x(415) & x(418) & x(428) & x(429) & x(430) & x(431) & x(432) & x(433) & x(436) & x(446) & x(457) & x(458) & x(459) & x(460) & x(461) & x(473) & x(474) & x(486) & x(487) & x(500) & x(501) & x(502) & x(515) & x(528) & x(529) & x(530) & x(555) & x(556) & x(557) & x(558) & x(584) & x(585) & x(612) & x(613) & x(619) & x(638) & x(640) & x(653) & x(679) & x(690) & x(691) & x(692) & x(693) & x(694) & x(695) & x(696) & x(706) & x(707) & x(708) & x(709) & x(721) & x(722) & x(723) & x(735) & x(736) & x(737) & x(739) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(764) & x(765) & x(766) & x(769) & x(770) & x(771) & x(772) & x(773) & x(774);
    y(174) <= not(p174_out);
    p174 : perceptron
        Generic map (
            WEIGHTS => "000000000000000000000000000000000010111110111111111111111111101100000000001110000000000001100010000000100000110011101111111111111111000000011110001111111111111111111",
            SHIFT => 3,
            B => 111,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p174_in,
            y(0) => p174_out,
            y(1 to 16 - 1) => dummy174
        );


    p175_in <= x(0) & x(2) & x(3) & x(4) & x(5) & x(11) & x(22) & x(23) & x(24) & x(27) & x(52) & x(54) & x(58) & x(75) & x(82) & x(84) & x(85) & x(110) & x(112) & x(139) & x(157) & x(159) & x(160) & x(196) & x(198) & x(199) & x(200) & x(201) & x(226) & x(227) & x(243) & x(249) & x(250) & x(254) & x(255) & x(266) & x(267) & x(268) & x(269) & x(270) & x(271) & x(277) & x(283) & x(284) & x(294) & x(295) & x(296) & x(309) & x(310) & x(312) & x(317) & x(318) & x(319) & x(320) & x(338) & x(339) & x(345) & x(347) & x(348) & x(353) & x(362) & x(364) & x(366) & x(367) & x(372) & x(373) & x(375) & x(380) & x(381) & x(382) & x(392) & x(402) & x(403) & x(404) & x(409) & x(416) & x(420) & x(430) & x(432) & x(433) & x(436) & x(437) & x(459) & x(460) & x(461) & x(487) & x(488) & x(508) & x(509) & x(514) & x(544) & x(571) & x(615) & x(616) & x(643) & x(644) & x(673) & x(675) & x(676) & x(677) & x(678) & x(679) & x(693) & x(694) & x(696) & x(699) & x(702) & x(705) & x(706) & x(707) & x(708) & x(709) & x(720) & x(721) & x(735) & x(736) & x(741) & x(742) & x(743) & x(744) & x(748) & x(754) & x(755) & x(758) & x(760) & x(764) & x(765) & x(766) & x(769) & x(770) & x(771) & x(773) & x(774) & x(779) & x(780) & x(781) & x(782) & x(783);
    y(175) <= not(p175_out);
    p175 : perceptron
        Generic map (
            WEIGHTS => "111111111111111111110001000000000000000000000000001111001111010011111111111011111111111001001111100000111110000011000000111110000000011111",
            SHIFT => 4,
            B => -8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p175_in,
            y(0) => p175_out,
            y(1 to 17 - 1) => dummy175
        );


    p176_in <= x(108) & x(191) & x(192) & x(193) & x(209) & x(210) & x(211) & x(212) & x(219) & x(220) & x(237) & x(238) & x(239) & x(247) & x(248) & x(266) & x(267) & x(276) & x(294) & x(295) & x(302) & x(322) & x(323) & x(328) & x(329) & x(330) & x(331) & x(332) & x(350) & x(378) & x(695) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(739) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(748) & x(749);
    y(176) <= not(p176_out);
    p176 : perceptron
        Generic map (
            WEIGHTS => "0111000011000110010000000000000000000000000000000",
            SHIFT => 4,
            B => -349,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p176_in,
            y(0) => p176_out,
            y(1 to 15 - 1) => dummy176
        );


    p177_in <= x(40) & x(43) & x(69) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(104) & x(105) & x(106) & x(107) & x(165) & x(192) & x(198) & x(216) & x(221) & x(222) & x(226) & x(248) & x(249) & x(250) & x(254) & x(268) & x(269) & x(277) & x(278) & x(282) & x(283) & x(295) & x(309) & x(310) & x(311) & x(312) & x(317) & x(318) & x(330) & x(331) & x(338) & x(339) & x(345) & x(348) & x(349) & x(350) & x(353) & x(354) & x(355) & x(358) & x(359) & x(362) & x(366) & x(377) & x(378) & x(379) & x(381) & x(382) & x(385) & x(386) & x(387) & x(390) & x(405) & x(406) & x(414) & x(418) & x(432) & x(433) & x(434) & x(435) & x(446) & x(460) & x(472) & x(473) & x(474) & x(484) & x(487) & x(488) & x(500) & x(501) & x(502) & x(509) & x(515) & x(528) & x(529) & x(530) & x(536) & x(537) & x(538) & x(553) & x(555) & x(556) & x(557) & x(558) & x(564) & x(566) & x(581) & x(583) & x(584) & x(585) & x(586) & x(591) & x(597) & x(598) & x(608) & x(611) & x(612) & x(619) & x(625) & x(638) & x(640) & x(651) & x(690) & x(691) & x(692) & x(693) & x(694) & x(695) & x(696) & x(706) & x(707) & x(708) & x(709) & x(710) & x(711) & x(712) & x(719) & x(720) & x(721) & x(722) & x(723) & x(735) & x(736) & x(737) & x(739) & x(741) & x(742) & x(743) & x(744) & x(748) & x(761) & x(764) & x(765) & x(766) & x(769) & x(770) & x(771) & x(772) & x(773) & x(774);
    y(177) <= not(p177_out);
    p177 : perceptron
        Generic map (
            WEIGHTS => "1111111111111110000000000000000000000111100111111111001111111101110111101000111000010000000000000000000000000000011111110000000111110000000010000000000",
            SHIFT => 4,
            B => -527,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p177_in,
            y(0) => p177_out,
            y(1 to 17 - 1) => dummy177
        );


    p178_in <= x(34) & x(35) & x(36) & x(37) & x(38) & x(39) & x(40) & x(41) & x(43) & x(47) & x(48) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(78) & x(79) & x(105) & x(118) & x(146) & x(171) & x(172) & x(173) & x(174) & x(197) & x(199) & x(200) & x(201) & x(202) & x(211) & x(228) & x(229) & x(248) & x(256) & x(268) & x(269) & x(276) & x(291) & x(295) & x(296) & x(297) & x(304) & x(310) & x(311) & x(315) & x(318) & x(323) & x(324) & x(342) & x(387) & x(388) & x(422) & x(437) & x(444) & x(446) & x(473) & x(474) & x(475) & x(479) & x(487) & x(501) & x(502) & x(507) & x(514) & x(515) & x(528) & x(529) & x(530) & x(535) & x(541) & x(542) & x(543) & x(556) & x(557) & x(558) & x(563) & x(570) & x(584) & x(591) & x(618) & x(619) & x(692) & x(693) & x(694) & x(695) & x(708) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(747) & x(748) & x(749) & x(769) & x(770) & x(771) & x(773);
    y(178) <= not(p178_out);
    p178 : perceptron
        Generic map (
            WEIGHTS => "111111111111111111111111111000000000001001000110001001100111001000001000110000111000010000111101111111110000",
            SHIFT => 4,
            B => 126,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p178_in,
            y(0) => p178_out,
            y(1 to 16 - 1) => dummy178
        );


    p179_in <= x(39) & x(44) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(78) & x(79) & x(90) & x(91) & x(93) & x(94) & x(95) & x(96) & x(104) & x(105) & x(108) & x(133) & x(181) & x(182) & x(183) & x(184) & x(192) & x(193) & x(194) & x(207) & x(208) & x(209) & x(213) & x(220) & x(221) & x(222) & x(248) & x(249) & x(276) & x(277) & x(305) & x(306) & x(323) & x(328) & x(329) & x(330) & x(331) & x(332) & x(341) & x(349) & x(359) & x(371) & x(372) & x(398) & x(399) & x(400) & x(401) & x(423) & x(427) & x(428) & x(429) & x(445) & x(472) & x(473) & x(479) & x(501) & x(502) & x(528) & x(529) & x(530) & x(535) & x(556) & x(557) & x(584) & x(611) & x(612) & x(638) & x(652) & x(654) & x(655) & x(656) & x(657) & x(681) & x(682) & x(683) & x(691) & x(692) & x(693) & x(694) & x(695) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(746) & x(747) & x(748) & x(749);
    y(179) <= not(p179_out);
    p179 : perceptron
        Generic map (
            WEIGHTS => "00000000000000000000011000000000000000000001111111011111110111000000000000000000000000111111111111111",
            SHIFT => 4,
            B => -326,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p179_in,
            y(0) => p179_out,
            y(1 to 16 - 1) => dummy179
        );


    p180_in <= x(34) & x(35) & x(36) & x(37) & x(38) & x(39) & x(40) & x(41) & x(42) & x(43) & x(44) & x(45) & x(46) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(79) & x(95) & x(96) & x(97) & x(98) & x(99) & x(100) & x(101) & x(102) & x(103) & x(104) & x(105) & x(106) & x(107) & x(108) & x(135) & x(136) & x(162) & x(163) & x(164) & x(165) & x(191) & x(192) & x(193) & x(194) & x(195) & x(219) & x(220) & x(221) & x(222) & x(247) & x(248) & x(249) & x(250) & x(276) & x(277) & x(302) & x(303) & x(304) & x(305) & x(328) & x(329) & x(330) & x(331) & x(332) & x(357) & x(358) & x(359) & x(360) & x(368) & x(369) & x(385) & x(386) & x(387) & x(388) & x(396) & x(414) & x(415) & x(416) & x(418) & x(443) & x(444) & x(446) & x(475) & x(487) & x(513) & x(514) & x(515) & x(516) & x(528) & x(530) & x(534) & x(541) & x(542) & x(543) & x(544) & x(571) & x(693) & x(694) & x(719) & x(721) & x(748) & x(749) & x(765);
    y(180) <= not(p180_out);
    p180 : perceptron
        Generic map (
            WEIGHTS => "000000000000000000000000000000000000000000000111111111111111111111000100000000011000010001001100000110000001111111",
            SHIFT => 4,
            B => -413,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p180_in,
            y(0) => p180_out,
            y(1 to 16 - 1) => dummy180
        );


    p181_in <= x(64) & x(78) & x(79) & x(104) & x(105) & x(138) & x(165) & x(166) & x(182) & x(183) & x(184) & x(193) & x(194) & x(210) & x(220) & x(221) & x(222) & x(247) & x(248) & x(249) & x(250) & x(275) & x(276) & x(277) & x(278) & x(303) & x(304) & x(305) & x(306) & x(307) & x(311) & x(321) & x(322) & x(333) & x(334) & x(340) & x(341) & x(348) & x(349) & x(350) & x(358) & x(359) & x(360) & x(361) & x(362) & x(376) & x(377) & x(378) & x(386) & x(387) & x(388) & x(390) & x(391) & x(405) & x(406) & x(418) & x(446) & x(454) & x(455) & x(501) & x(529) & x(530) & x(557) & x(558) & x(584) & x(585) & x(612) & x(657) & x(692) & x(695) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(724) & x(746) & x(747) & x(748) & x(749);
    y(181) <= not(p181_out);
    p181 : perceptron
        Generic map (
            WEIGHTS => "1111100000000000000000000000001000000000111000001110000001111111111000000000000000",
            SHIFT => 4,
            B => -466,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p181_in,
            y(0) => p181_out,
            y(1 to 16 - 1) => dummy181
        );


    p182_in <= x(67) & x(68) & x(69) & x(70) & x(72) & x(73) & x(76) & x(77) & x(78) & x(79) & x(80) & x(94) & x(96) & x(101) & x(102) & x(103) & x(104) & x(105) & x(106) & x(121) & x(147) & x(148) & x(192) & x(219) & x(220) & x(247) & x(248) & x(249) & x(250) & x(275) & x(276) & x(277) & x(287) & x(288) & x(289) & x(290) & x(291) & x(294) & x(303) & x(304) & x(307) & x(315) & x(316) & x(317) & x(320) & x(327) & x(328) & x(334) & x(338) & x(339) & x(346) & x(347) & x(349) & x(353) & x(354) & x(355) & x(362) & x(366) & x(394) & x(397) & x(436) & x(463) & x(468) & x(469) & x(473) & x(474) & x(498) & x(501) & x(502) & x(508) & x(525) & x(526) & x(528) & x(529) & x(530) & x(536) & x(537) & x(538) & x(553) & x(557) & x(558) & x(564) & x(565) & x(581) & x(584) & x(592) & x(593) & x(594) & x(612) & x(621) & x(649) & x(656) & x(657) & x(660) & x(674) & x(688) & x(739) & x(742) & x(744) & x(745) & x(746) & x(770) & x(773) & x(774);
    y(182) <= not(p182_out);
    p182 : perceptron
        Generic map (
            WEIGHTS => "00000000000000000000001111111111111110111111111100111111100111000000000000000000000000000001111100000000",
            SHIFT => 4,
            B => -550,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p182_in,
            y(0) => p182_out,
            y(1 to 16 - 1) => dummy182
        );


    p183_in <= x(35) & x(37) & x(40) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(90) & x(91) & x(92) & x(93) & x(94) & x(108) & x(109) & x(165) & x(166) & x(171) & x(172) & x(188) & x(192) & x(193) & x(194) & x(199) & x(200) & x(219) & x(220) & x(221) & x(222) & x(247) & x(248) & x(249) & x(250) & x(275) & x(276) & x(277) & x(295) & x(296) & x(297) & x(298) & x(299) & x(300) & x(301) & x(320) & x(325) & x(326) & x(327) & x(328) & x(331) & x(332) & x(348) & x(350) & x(404) & x(446) & x(450) & x(474) & x(475) & x(535) & x(706) & x(707) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(735) & x(744) & x(745) & x(746) & x(747) & x(748);
    y(183) <= not(p183_out);
    p183 : perceptron
        Generic map (
            WEIGHTS => "11111111111111100110011110011111111111000000010000001110000000000000000000",
            SHIFT => 4,
            B => 42,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p183_in,
            y(0) => p183_out,
            y(1 to 16 - 1) => dummy183
        );


    p184_in <= x(39) & x(40) & x(45) & x(49) & x(63) & x(64) & x(66) & x(68) & x(95) & x(96) & x(100) & x(103) & x(108) & x(163) & x(165) & x(192) & x(194) & x(220) & x(221) & x(222) & x(242) & x(248) & x(249) & x(250) & x(268) & x(269) & x(270) & x(276) & x(277) & x(278) & x(297) & x(298) & x(299) & x(300) & x(301) & x(302) & x(303) & x(305) & x(309) & x(323) & x(325) & x(326) & x(327) & x(328) & x(329) & x(330) & x(331) & x(332) & x(350) & x(357) & x(358) & x(359) & x(360) & x(394) & x(400) & x(446) & x(455) & x(456) & x(457) & x(458) & x(459) & x(475) & x(483) & x(511) & x(512) & x(514) & x(535) & x(540) & x(541) & x(542) & x(543) & x(552) & x(570) & x(571) & x(572) & x(656) & x(657) & x(658) & x(659) & x(660) & x(682) & x(683) & x(684) & x(685) & x(686) & x(687) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(740) & x(742) & x(744) & x(745) & x(746);
    y(184) <= not(p184_out);
    p184 : perceptron
        Generic map (
            WEIGHTS => "0000000000001000000010001110001111111011111111111111110100000100010000000001111111111111111111111",
            SHIFT => 3,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p184_in,
            y(0) => p184_out,
            y(1 to 15 - 1) => dummy184
        );


    p185_in <= x(35) & x(39) & x(40) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(75) & x(91) & x(92) & x(93) & x(94) & x(95) & x(126) & x(131) & x(135) & x(136) & x(164) & x(165) & x(171) & x(172) & x(173) & x(192) & x(193) & x(197) & x(199) & x(200) & x(201) & x(202) & x(220) & x(221) & x(227) & x(228) & x(229) & x(232) & x(238) & x(245) & x(248) & x(249) & x(250) & x(254) & x(255) & x(266) & x(269) & x(270) & x(271) & x(274) & x(276) & x(277) & x(278) & x(283) & x(305) & x(307) & x(320) & x(333) & x(334) & x(347) & x(348) & x(349) & x(358) & x(361) & x(362) & x(381) & x(409) & x(423) & x(450) & x(457) & x(458) & x(473) & x(474) & x(478) & x(501) & x(502) & x(506) & x(507) & x(511) & x(516) & x(526) & x(529) & x(534) & x(535) & x(543) & x(545) & x(557) & x(573) & x(574) & x(582) & x(584) & x(611) & x(612) & x(638) & x(647) & x(648) & x(656) & x(657) & x(660) & x(675) & x(676) & x(677) & x(679) & x(680) & x(697) & x(706) & x(707) & x(708) & x(718) & x(734) & x(735) & x(736) & x(737) & x(769) & x(770) & x(773);
    y(185) <= not(p185_out);
    p185 : perceptron
        Generic map (
            WEIGHTS => "0000000000000000000011111111111111111111011111101111111111111111011111100001001100001100000000001111111111011101111111",
            SHIFT => 4,
            B => 485,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p185_in,
            y(0) => p185_out,
            y(1 to 17 - 1) => dummy185
        );


    p186_in <= x(44) & x(64) & x(66) & x(67) & x(68) & x(70) & x(91) & x(92) & x(93) & x(94) & x(95) & x(96) & x(98) & x(99) & x(100) & x(101) & x(106) & x(107) & x(108) & x(151) & x(178) & x(179) & x(184) & x(193) & x(194) & x(198) & x(199) & x(221) & x(222) & x(226) & x(227) & x(228) & x(248) & x(249) & x(250) & x(276) & x(277) & x(278) & x(298) & x(302) & x(305) & x(306) & x(309) & x(314) & x(322) & x(323) & x(324) & x(325) & x(326) & x(327) & x(328) & x(329) & x(330) & x(331) & x(348) & x(350) & x(357) & x(375) & x(379) & x(382) & x(390) & x(394) & x(403) & x(406) & x(409) & x(418) & x(430) & x(431) & x(435) & x(446) & x(462) & x(472) & x(473) & x(474) & x(490) & x(495) & x(497) & x(500) & x(501) & x(502) & x(509) & x(523) & x(528) & x(529) & x(536) & x(537) & x(539) & x(540) & x(543) & x(548) & x(549) & x(550) & x(552) & x(553) & x(556) & x(557) & x(558) & x(564) & x(565) & x(569) & x(571) & x(579) & x(583) & x(584) & x(585) & x(600) & x(610) & x(611) & x(612) & x(622) & x(624) & x(636) & x(637) & x(638) & x(639) & x(649) & x(650) & x(651) & x(691) & x(692) & x(693) & x(695) & x(697) & x(706) & x(707) & x(708) & x(714) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(735) & x(736) & x(737) & x(738) & x(739) & x(740) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(765) & x(769) & x(770) & x(771) & x(773);
    y(186) <= not(p186_out);
    p186 : perceptron
        Generic map (
            WEIGHTS => "00000000000000001110000001100111000000110011111111111101101101011000101000100000000000000000000000000000000000000000001111011111111111111111111111111111",
            SHIFT => 3,
            B => -213,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p186_in,
            y(0) => p186_out,
            y(1 to 16 - 1) => dummy186
        );


    p187_in <= x(63) & x(64) & x(104) & x(105) & x(177) & x(191) & x(192) & x(198) & x(219) & x(221) & x(226) & x(227) & x(248) & x(249) & x(254) & x(265) & x(266) & x(267) & x(270) & x(276) & x(277) & x(293) & x(294) & x(295) & x(298) & x(303) & x(309) & x(310) & x(320) & x(328) & x(329) & x(338) & x(339) & x(348) & x(349) & x(350) & x(351) & x(361) & x(362) & x(366) & x(376) & x(377) & x(378) & x(379) & x(381) & x(385) & x(386) & x(403) & x(404) & x(405) & x(414) & x(418) & x(432) & x(433) & x(446) & x(455) & x(460) & x(461) & x(464) & x(474) & x(484) & x(535) & x(543) & x(544) & x(545) & x(572) & x(595) & x(623) & x(632) & x(633) & x(634) & x(647) & x(652) & x(655) & x(656) & x(657) & x(664) & x(737) & x(739) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(764) & x(765) & x(769) & x(770) & x(773) & x(774);
    y(187) <= not(p187_out);
    p187 : perceptron
        Generic map (
            WEIGHTS => "1111111011001100000110000000100001111000111110011100110011100100001111111111100000000000000",
            SHIFT => 4,
            B => -138,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p187_in,
            y(0) => p187_out,
            y(1 to 16 - 1) => dummy187
        );


    p188_in <= x(69) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(100) & x(101) & x(102) & x(103) & x(104) & x(105) & x(106) & x(107) & x(108) & x(121) & x(162) & x(163) & x(164) & x(165) & x(188) & x(189) & x(191) & x(192) & x(193) & x(194) & x(195) & x(201) & x(204) & x(210) & x(211) & x(217) & x(220) & x(221) & x(222) & x(242) & x(243) & x(244) & x(245) & x(248) & x(249) & x(250) & x(269) & x(276) & x(277) & x(278) & x(283) & x(303) & x(305) & x(330) & x(331) & x(332) & x(341) & x(342) & x(356) & x(357) & x(359) & x(370) & x(390) & x(398) & x(403) & x(418) & x(431) & x(438) & x(446) & x(450) & x(466) & x(467) & x(472) & x(473) & x(474) & x(479) & x(486) & x(487) & x(501) & x(502) & x(507) & x(513) & x(514) & x(515) & x(516) & x(528) & x(529) & x(535) & x(536) & x(556) & x(557) & x(563) & x(564) & x(584) & x(591) & x(592) & x(619) & x(620) & x(636) & x(647) & x(648) & x(649) & x(677) & x(690) & x(691) & x(692) & x(693) & x(694) & x(695) & x(708) & x(718) & x(719) & x(720) & x(721) & x(722) & x(746) & x(764) & x(765) & x(766) & x(769) & x(770);
    y(188) <= not(p188_out);
    p188 : perceptron
        Generic map (
            WEIGHTS => "111111111111111111000000000000001100000000000000001011100111000101000000000110001111000000000000000000111111011111100000",
            SHIFT => 4,
            B => -420,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p188_in,
            y(0) => p188_out,
            y(1 to 17 - 1) => dummy188
        );


    p189_in <= x(79) & x(102) & x(105) & x(146) & x(163) & x(172) & x(173) & x(174) & x(182) & x(183) & x(184) & x(197) & x(202) & x(209) & x(210) & x(211) & x(212) & x(228) & x(229) & x(237) & x(238) & x(239) & x(240) & x(248) & x(250) & x(256) & x(275) & x(276) & x(283) & x(289) & x(291) & x(303) & x(304) & x(310) & x(311) & x(312) & x(315) & x(331) & x(339) & x(341) & x(342) & x(343) & x(349) & x(350) & x(359) & x(369) & x(437) & x(450) & x(473) & x(479) & x(501) & x(502) & x(507) & x(528) & x(529) & x(530) & x(535) & x(556) & x(557) & x(558) & x(563) & x(584) & x(591) & x(612) & x(619) & x(620) & x(676) & x(690) & x(691) & x(692) & x(693) & x(694) & x(695) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(724) & x(735) & x(736) & x(745) & x(746) & x(747) & x(748) & x(749) & x(762) & x(764) & x(766) & x(767) & x(768) & x(769) & x(770) & x(771) & x(772) & x(773) & x(774);
    y(189) <= not(p189_out);
    p189 : perceptron
        Generic map (
            WEIGHTS => "0000000011100111100111111011011110001101111111000000000000000000000111111111111111001111100000000000",
            SHIFT => 4,
            B => -321,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p189_in,
            y(0) => p189_out,
            y(1 to 16 - 1) => dummy189
        );


    p190_in <= x(124) & x(125) & x(151) & x(152) & x(163) & x(181) & x(182) & x(190) & x(192) & x(209) & x(210) & x(211) & x(212) & x(213) & x(220) & x(233) & x(239) & x(240) & x(248) & x(249) & x(260) & x(277) & x(284) & x(287) & x(305) & x(320) & x(321) & x(333) & x(334) & x(340) & x(359) & x(361) & x(362) & x(387) & x(401) & x(427) & x(428) & x(429) & x(430) & x(453) & x(455) & x(462) & x(463) & x(479) & x(481) & x(482) & x(483) & x(489) & x(490) & x(501) & x(507) & x(517) & x(528) & x(529) & x(557) & x(584) & x(706) & x(707) & x(708) & x(734) & x(736) & x(737) & x(738) & x(739) & x(740) & x(742) & x(743) & x(770);
    y(190) <= not(p190_out);
    p190 : perceptron
        Generic map (
            WEIGHTS => "00001001100000110011111111111101100000000111000110110000111111111111",
            SHIFT => 4,
            B => 245,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p190_in,
            y(0) => p190_out,
            y(1 to 16 - 1) => dummy190
        );


    p191_in <= x(105) & x(106) & x(193) & x(198) & x(220) & x(221) & x(247) & x(248) & x(249) & x(250) & x(264) & x(275) & x(276) & x(277) & x(303) & x(304) & x(305) & x(306) & x(307) & x(309) & x(310) & x(311) & x(320) & x(321) & x(322) & x(332) & x(333) & x(334) & x(338) & x(339) & x(347) & x(348) & x(349) & x(350) & x(351) & x(361) & x(362) & x(366) & x(375) & x(376) & x(377) & x(378) & x(394) & x(433) & x(444) & x(450) & x(473) & x(501) & x(506) & x(507) & x(528) & x(529) & x(530) & x(534) & x(535) & x(556) & x(557) & x(563) & x(584) & x(591) & x(638) & x(647) & x(655) & x(656) & x(657) & x(658) & x(674) & x(675) & x(693) & x(695) & x(708) & x(721) & x(722) & x(723) & x(735) & x(736) & x(737) & x(738) & x(739) & x(742) & x(743) & x(744) & x(745) & x(746) & x(765) & x(769) & x(770) & x(772) & x(773) & x(774);
    y(191) <= not(p191_out);
    p191 : perceptron
        Generic map (
            WEIGHTS => "001011111101111111100011111100111111101111011100110001100101011111111101110000000000000000",
            SHIFT => 4,
            B => 84,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p191_in,
            y(0) => p191_out,
            y(1 to 16 - 1) => dummy191
        );


    p192_in <= x(69) & x(71) & x(166) & x(192) & x(193) & x(194) & x(220) & x(221) & x(222) & x(247) & x(248) & x(249) & x(250) & x(275) & x(276) & x(277) & x(278) & x(305) & x(306) & x(320) & x(321) & x(333) & x(334) & x(347) & x(348) & x(349) & x(350) & x(351) & x(366) & x(375) & x(376) & x(377) & x(378) & x(404) & x(405) & x(406) & x(453) & x(455) & x(473) & x(474) & x(501) & x(502) & x(507) & x(529) & x(557) & x(558) & x(584) & x(612) & x(638) & x(656) & x(657) & x(692) & x(693) & x(694) & x(695) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(747) & x(748) & x(749);
    y(192) <= not(p192_out);
    p192 : perceptron
        Generic map (
            WEIGHTS => "1111111111111111111111111111011111110000001000000111111111111111",
            SHIFT => 4,
            B => 484,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p192_in,
            y(0) => p192_out,
            y(1 to 16 - 1) => dummy192
        );


    p193_in <= x(35) & x(37) & x(38) & x(39) & x(40) & x(41) & x(45) & x(46) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(79) & x(98) & x(99) & x(100) & x(101) & x(102) & x(103) & x(104) & x(105) & x(106) & x(107) & x(108) & x(155) & x(157) & x(198) & x(226) & x(258) & x(280) & x(284) & x(307) & x(309) & x(310) & x(311) & x(312) & x(333) & x(337) & x(338) & x(339) & x(361) & x(362) & x(366) & x(375) & x(380) & x(388) & x(390) & x(394) & x(401) & x(403) & x(410) & x(414) & x(416) & x(418) & x(429) & x(446) & x(450) & x(473) & x(474) & x(475) & x(489) & x(501) & x(502) & x(506) & x(507) & x(519) & x(528) & x(529) & x(530) & x(534) & x(535) & x(555) & x(556) & x(557) & x(584) & x(591) & x(619) & x(647) & x(648) & x(674) & x(675) & x(676) & x(677) & x(678) & x(693) & x(694) & x(695) & x(705) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(732) & x(747) & x(748) & x(749) & x(764) & x(765) & x(769) & x(770) & x(773) & x(774);
    y(193) <= not(p193_out);
    p193 : perceptron
        Generic map (
            WEIGHTS => "0000000000000000000000000000000000000111111111111111111100011000001010111111001111001111000000000000000000000000111111",
            SHIFT => 5,
            B => -842,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p193_in,
            y(0) => p193_out,
            y(1 to 18 - 1) => dummy193
        );


    p194_in <= x(35) & x(63) & x(64) & x(67) & x(108) & x(163) & x(171) & x(191) & x(192) & x(197) & x(210) & x(211) & x(238) & x(239) & x(277) & x(289) & x(290) & x(305) & x(329) & x(331) & x(333) & x(334) & x(338) & x(349) & x(400) & x(425) & x(435) & x(450) & x(488) & x(507) & x(516) & x(535) & x(563) & x(591) & x(647) & x(675) & x(703) & x(709) & x(713) & x(715) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(732) & x(733) & x(734) & x(736) & x(737) & x(738) & x(739) & x(740) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(748) & x(749) & x(770);
    y(194) <= not(p194_out);
    p194 : perceptron
        Generic map (
            WEIGHTS => "000001111100001001001101111111111111100000000000000000000000000000",
            SHIFT => 5,
            B => -397,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p194_in,
            y(0) => p194_out,
            y(1 to 17 - 1) => dummy194
        );


    p195_in <= x(35) & x(37) & x(38) & x(39) & x(40) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(79) & x(90) & x(91) & x(92) & x(93) & x(94) & x(136) & x(181) & x(182) & x(183) & x(184) & x(210) & x(211) & x(249) & x(277) & x(294) & x(297) & x(298) & x(299) & x(300) & x(302) & x(303) & x(307) & x(325) & x(326) & x(327) & x(329) & x(330) & x(331) & x(332) & x(350) & x(355) & x(361) & x(369) & x(371) & x(378) & x(396) & x(397) & x(424) & x(425) & x(436) & x(437) & x(464) & x(529) & x(556) & x(557) & x(584) & x(596) & x(597) & x(611) & x(612) & x(624) & x(625) & x(638) & x(690) & x(691) & x(692) & x(693) & x(695) & x(719);
    y(195) <= not(p195_out);
    p195 : perceptron
        Generic map (
            WEIGHTS => "11111111111111111111011111111100000000000000100001000000011111111111000000",
            SHIFT => 4,
            B => 144,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p195_in,
            y(0) => p195_out,
            y(1 to 16 - 1) => dummy195
        );


    p196_in <= x(44) & x(66) & x(67) & x(68) & x(69) & x(70) & x(91) & x(93) & x(94) & x(95) & x(96) & x(97) & x(133) & x(134) & x(135) & x(153) & x(154) & x(156) & x(166) & x(179) & x(180) & x(182) & x(183) & x(193) & x(198) & x(221) & x(248) & x(249) & x(250) & x(275) & x(276) & x(277) & x(278) & x(303) & x(304) & x(305) & x(306) & x(324) & x(333) & x(334) & x(342) & x(361) & x(362) & x(370) & x(371) & x(372) & x(373) & x(389) & x(390) & x(396) & x(397) & x(399) & x(401) & x(418) & x(421) & x(433) & x(445) & x(446) & x(450) & x(471) & x(473) & x(474) & x(479) & x(498) & x(500) & x(501) & x(502) & x(507) & x(528) & x(529) & x(535) & x(536) & x(541) & x(542) & x(556) & x(557) & x(558) & x(563) & x(564) & x(569) & x(579) & x(583) & x(584) & x(591) & x(596) & x(612) & x(619) & x(620) & x(625) & x(627) & x(640) & x(647) & x(670) & x(693) & x(694) & x(739) & x(777);
    y(196) <= not(p196_out);
    p196 : perceptron
        Generic map (
            WEIGHTS => "0000000000001110000000001000000000000100100111100111101000000000000000000000000000000000000011110",
            SHIFT => 4,
            B => -856,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p196_in,
            y(0) => p196_out,
            y(1 to 16 - 1) => dummy196
        );


    p197_in <= x(34) & x(35) & x(36) & x(37) & x(38) & x(39) & x(40) & x(41) & x(44) & x(45) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(79) & x(90) & x(91) & x(92) & x(93) & x(94) & x(95) & x(96) & x(104) & x(105) & x(106) & x(109) & x(165) & x(166) & x(171) & x(172) & x(191) & x(192) & x(193) & x(194) & x(199) & x(200) & x(210) & x(211) & x(219) & x(220) & x(221) & x(222) & x(247) & x(248) & x(249) & x(250) & x(267) & x(268) & x(275) & x(276) & x(277) & x(292) & x(294) & x(295) & x(296) & x(297) & x(298) & x(299) & x(300) & x(301) & x(302) & x(306) & x(320) & x(322) & x(323) & x(324) & x(325) & x(326) & x(327) & x(328) & x(348) & x(397) & x(418) & x(425) & x(445) & x(450) & x(507) & x(515) & x(516) & x(535) & x(542) & x(543) & x(544) & x(563) & x(591) & x(611) & x(619) & x(675) & x(676) & x(677) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(739) & x(742) & x(744) & x(745) & x(746) & x(747) & x(748);
    y(197) <= not(p197_out);
    p197 : perceptron
        Generic map (
            WEIGHTS => "00000000000000000000000000000000000000100110000111100000000110000111111111001111111011101100100011011111111111111111",
            SHIFT => 4,
            B => -387,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p197_in,
            y(0) => p197_out,
            y(1 to 16 - 1) => dummy197
        );


    p198_in <= x(0) & x(1) & x(2) & x(3) & x(4) & x(5) & x(6) & x(7) & x(8) & x(9) & x(10) & x(11) & x(12) & x(15) & x(16) & x(17) & x(18) & x(19) & x(20) & x(21) & x(22) & x(23) & x(24) & x(25) & x(26) & x(27) & x(28) & x(29) & x(30) & x(31) & x(32) & x(33) & x(44) & x(52) & x(53) & x(54) & x(55) & x(56) & x(57) & x(58) & x(59) & x(61) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(82) & x(83) & x(84) & x(85) & x(87) & x(88) & x(91) & x(92) & x(93) & x(94) & x(95) & x(96) & x(104) & x(105) & x(106) & x(110) & x(111) & x(112) & x(113) & x(115) & x(139) & x(140) & x(141) & x(142) & x(167) & x(168) & x(169) & x(192) & x(193) & x(194) & x(196) & x(220) & x(221) & x(222) & x(248) & x(249) & x(250) & x(276) & x(277) & x(278) & x(283) & x(302) & x(305) & x(306) & x(310) & x(311) & x(330) & x(331) & x(338) & x(339) & x(358) & x(359) & x(364) & x(370) & x(386) & x(390) & x(392) & x(396) & x(397) & x(414) & x(419) & x(420) & x(445) & x(448) & x(449) & x(473) & x(474) & x(476) & x(479) & x(501) & x(502) & x(503) & x(504) & x(507) & x(528) & x(529) & x(532) & x(535) & x(557) & x(560) & x(563) & x(584) & x(587) & x(588) & x(591) & x(615) & x(616) & x(617) & x(619) & x(643) & x(644) & x(645) & x(671) & x(672) & x(673) & x(691) & x(692) & x(694) & x(698) & x(699) & x(700) & x(701) & x(702) & x(707) & x(708) & x(709) & x(710) & x(711) & x(712) & x(725) & x(726) & x(727) & x(728) & x(729) & x(730) & x(731) & x(735) & x(736) & x(737) & x(738) & x(739) & x(740) & x(752) & x(753) & x(754) & x(755) & x(756) & x(757) & x(758) & x(759) & x(760) & x(767) & x(768) & x(769) & x(770) & x(771) & x(772) & x(779) & x(780) & x(781) & x(782) & x(783);
    y(198) <= not(p198_out);
    p198 : perceptron
        Generic map (
            WEIGHTS => "11111111111111111111111111111111011111111100000000001111110000000001111111111110001000000000010000110011111011111101100100011000100100110111011111111111111000000111111100000011111111100000011111",
            SHIFT => 5,
            B => 1586,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p198_in,
            y(0) => p198_out,
            y(1 to 18 - 1) => dummy198
        );


    p199_in <= x(35) & x(39) & x(40) & x(44) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(70) & x(78) & x(79) & x(90) & x(91) & x(92) & x(93) & x(94) & x(95) & x(96) & x(104) & x(105) & x(106) & x(152) & x(171) & x(179) & x(180) & x(184) & x(199) & x(200) & x(226) & x(227) & x(228) & x(248) & x(249) & x(254) & x(255) & x(266) & x(267) & x(276) & x(294) & x(295) & x(296) & x(297) & x(311) & x(312) & x(322) & x(323) & x(347) & x(348) & x(349) & x(361) & x(366) & x(371) & x(375) & x(376) & x(399) & x(400) & x(403) & x(405) & x(426) & x(427) & x(428) & x(431) & x(432) & x(433) & x(455) & x(456) & x(457) & x(459) & x(460) & x(473) & x(487) & x(488) & x(501) & x(502) & x(514) & x(515) & x(529) & x(535) & x(542) & x(557) & x(584) & x(607) & x(623) & x(626) & x(627) & x(653) & x(655) & x(656) & x(657) & x(667) & x(675) & x(676) & x(677) & x(678) & x(690) & x(695) & x(705) & x(706) & x(707) & x(708) & x(718) & x(719) & x(720) & x(721) & x(722) & x(732) & x(735) & x(737) & x(748) & x(749) & x(770) & x(773);
    y(199) <= not(p199_out);
    p199 : perceptron
        Generic map (
            WEIGHTS => "0000000000000000000000000100011111001111011111111000111001100111000111000000000010000000000001111001111000000110011",
            SHIFT => 4,
            B => -262,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p199_in,
            y(0) => p199_out,
            y(1 to 16 - 1) => dummy199
        );


    p200_in <= x(0) & x(1) & x(2) & x(3) & x(4) & x(5) & x(6) & x(7) & x(8) & x(9) & x(10) & x(11) & x(12) & x(15) & x(16) & x(17) & x(18) & x(19) & x(20) & x(21) & x(22) & x(23) & x(24) & x(25) & x(26) & x(27) & x(28) & x(29) & x(30) & x(31) & x(32) & x(33) & x(34) & x(35) & x(36) & x(37) & x(38) & x(39) & x(40) & x(41) & x(45) & x(46) & x(49) & x(52) & x(53) & x(54) & x(55) & x(56) & x(57) & x(58) & x(59) & x(61) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(82) & x(83) & x(84) & x(85) & x(87) & x(88) & x(92) & x(99) & x(110) & x(111) & x(112) & x(113) & x(115) & x(123) & x(124) & x(131) & x(132) & x(139) & x(140) & x(141) & x(142) & x(147) & x(148) & x(149) & x(150) & x(165) & x(167) & x(168) & x(169) & x(196) & x(221) & x(222) & x(227) & x(248) & x(249) & x(250) & x(254) & x(266) & x(276) & x(277) & x(293) & x(294) & x(297) & x(301) & x(302) & x(303) & x(326) & x(327) & x(329) & x(330) & x(331) & x(332) & x(342) & x(353) & x(361) & x(364) & x(381) & x(385) & x(386) & x(387) & x(392) & x(404) & x(409) & x(410) & x(413) & x(414) & x(415) & x(416) & x(419) & x(420) & x(425) & x(432) & x(433) & x(434) & x(436) & x(443) & x(444) & x(446) & x(448) & x(449) & x(453) & x(460) & x(463) & x(464) & x(469) & x(473) & x(474) & x(475) & x(476) & x(485) & x(488) & x(491) & x(492) & x(495) & x(501) & x(502) & x(503) & x(504) & x(514) & x(528) & x(529) & x(530) & x(531) & x(532) & x(542) & x(543) & x(544) & x(557) & x(558) & x(560) & x(571) & x(572) & x(573) & x(580) & x(582) & x(583) & x(584) & x(587) & x(588) & x(601) & x(602) & x(603) & x(607) & x(609) & x(610) & x(611) & x(612) & x(615) & x(616) & x(617) & x(638) & x(639) & x(643) & x(644) & x(645) & x(653) & x(665) & x(666) & x(671) & x(672) & x(673) & x(675) & x(676) & x(677) & x(678) & x(691) & x(692) & x(698) & x(699) & x(700) & x(701) & x(702) & x(705) & x(708) & x(709) & x(712) & x(721) & x(725) & x(726) & x(727) & x(728) & x(729) & x(730) & x(731) & x(736) & x(738) & x(739) & x(740) & x(741) & x(742) & x(743) & x(744) & x(752) & x(753) & x(754) & x(755) & x(756) & x(757) & x(758) & x(759) & x(760) & x(779) & x(780) & x(781) & x(782) & x(783);
    y(200) <= not(p200_out);
    p200 : perceptron
        Generic map (
            WEIGHTS => "1111111111111111111111111111111100000000000111111111000000000000000111111001111111001111111101111000000000000111111111101111000111100001111111001111111011111111011111111110001110001111110001111111111111011111000011111110000011111110000000011111111111111",
            SHIFT => 4,
            B => 165,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p200_in,
            y(0) => p200_out,
            y(1 to 18 - 1) => dummy200
        );


    p201_in <= x(74) & x(91) & x(93) & x(94) & x(95) & x(96) & x(166) & x(193) & x(205) & x(206) & x(220) & x(221) & x(248) & x(249) & x(250) & x(273) & x(274) & x(276) & x(277) & x(278) & x(301) & x(302) & x(305) & x(306) & x(332) & x(334) & x(339) & x(362) & x(367) & x(370) & x(371) & x(374) & x(385) & x(390) & x(398) & x(401) & x(411) & x(414) & x(415) & x(416) & x(418) & x(429) & x(445) & x(446) & x(457) & x(473) & x(474) & x(479) & x(500) & x(501) & x(502) & x(507) & x(528) & x(529) & x(530) & x(535) & x(537) & x(541) & x(555) & x(556) & x(557) & x(558) & x(567) & x(568) & x(569) & x(583) & x(584) & x(585) & x(591) & x(595) & x(610) & x(611) & x(612) & x(619) & x(627) & x(638) & x(640) & x(655) & x(656) & x(657) & x(658) & x(670) & x(692) & x(693) & x(694) & x(719) & x(721) & x(769) & x(771);
    y(201) <= not(p201_out);
    p201 : perceptron
        Generic map (
            WEIGHTS => "01111111111111111111111111111000010000001011011111111111111111111111111111111111100000011",
            SHIFT => 4,
            B => 853,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p201_in,
            y(0) => p201_out,
            y(1 to 16 - 1) => dummy201
        );


    p202_in <= x(37) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(90) & x(92) & x(105) & x(117) & x(118) & x(125) & x(145) & x(147) & x(148) & x(149) & x(152) & x(164) & x(165) & x(166) & x(171) & x(172) & x(173) & x(174) & x(175) & x(192) & x(193) & x(194) & x(198) & x(200) & x(220) & x(221) & x(222) & x(247) & x(248) & x(249) & x(250) & x(254) & x(264) & x(276) & x(277) & x(289) & x(291) & x(292) & x(295) & x(297) & x(298) & x(299) & x(300) & x(302) & x(303) & x(304) & x(315) & x(316) & x(317) & x(319) & x(320) & x(323) & x(326) & x(327) & x(330) & x(331) & x(332) & x(340) & x(341) & x(342) & x(343) & x(344) & x(347) & x(350) & x(357) & x(360) & x(361) & x(362) & x(368) & x(378) & x(386) & x(387) & x(394) & x(415) & x(416) & x(446) & x(450) & x(479) & x(490) & x(502) & x(507) & x(529) & x(534) & x(535) & x(557) & x(562) & x(563) & x(570) & x(584) & x(591) & x(598) & x(599) & x(612) & x(618) & x(619) & x(647) & x(648) & x(675) & x(707) & x(709) & x(710) & x(711) & x(712) & x(715) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(734) & x(735) & x(736) & x(737) & x(738) & x(739) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(769) & x(770);
    y(202) <= not(p202_out);
    p202 : perceptron
        Generic map (
            WEIGHTS => "000000000001111111100011111000010000000000000011111111000001111110000001011101000001111111111110110011111100000000000000000000000000",
            SHIFT => 4,
            B => -378,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p202_in,
            y(0) => p202_out,
            y(1 to 17 - 1) => dummy202
        );


    p203_in <= x(34) & x(35) & x(36) & x(37) & x(38) & x(39) & x(40) & x(41) & x(46) & x(47) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(79) & x(91) & x(96) & x(97) & x(98) & x(99) & x(100) & x(101) & x(102) & x(103) & x(104) & x(105) & x(106) & x(107) & x(108) & x(162) & x(163) & x(190) & x(191) & x(192) & x(193) & x(210) & x(211) & x(218) & x(219) & x(220) & x(221) & x(238) & x(247) & x(248) & x(249) & x(305) & x(330) & x(331) & x(334) & x(357) & x(358) & x(359) & x(386) & x(387) & x(415) & x(418) & x(425) & x(446) & x(474) & x(487) & x(501) & x(502) & x(514) & x(515) & x(516) & x(528) & x(529) & x(530) & x(535) & x(542) & x(543) & x(544) & x(556) & x(557) & x(558) & x(584) & x(586) & x(612) & x(693) & x(695) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(739) & x(740) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(748) & x(749);
    y(203) <= not(p203_out);
    p203 : perceptron
        Generic map (
            WEIGHTS => "0000000000000000000000000000000000000000001111110011110111100100000011110110001111000111111000000000000000000000",
            SHIFT => 4,
            B => -742,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p203_in,
            y(0) => p203_out,
            y(1 to 16 - 1) => dummy203
        );


    p204_in <= x(34) & x(35) & x(36) & x(37) & x(38) & x(39) & x(40) & x(41) & x(44) & x(45) & x(46) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(79) & x(90) & x(91) & x(94) & x(95) & x(96) & x(97) & x(98) & x(99) & x(100) & x(101) & x(102) & x(103) & x(104) & x(105) & x(106) & x(107) & x(108) & x(122) & x(124) & x(125) & x(126) & x(127) & x(152) & x(153) & x(154) & x(155) & x(162) & x(163) & x(164) & x(177) & x(179) & x(182) & x(183) & x(190) & x(191) & x(192) & x(193) & x(210) & x(211) & x(219) & x(236) & x(238) & x(241) & x(242) & x(243) & x(247) & x(248) & x(249) & x(263) & x(264) & x(269) & x(270) & x(294) & x(307) & x(322) & x(334) & x(345) & x(349) & x(358) & x(359) & x(360) & x(361) & x(362) & x(370) & x(373) & x(385) & x(387) & x(388) & x(397) & x(398) & x(399) & x(401) & x(418) & x(437) & x(446) & x(464) & x(488) & x(489) & x(492) & x(514) & x(515) & x(516) & x(523) & x(541) & x(542) & x(543) & x(544) & x(570) & x(571) & x(572) & x(591) & x(623) & x(690) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(732) & x(739) & x(741) & x(745) & x(746) & x(747) & x(748) & x(749);
    y(204) <= not(p204_out);
    p204 : perceptron
        Generic map (
            WEIGHTS => "000000000000000000000000000000000000000000000000000000011100001111001101111111111010110000111100011111111001000000000000010000000000000000",
            SHIFT => 3,
            B => -532,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p204_in,
            y(0) => p204_out,
            y(1 to 16 - 1) => dummy204
        );


    p205_in <= x(165) & x(192) & x(221) & x(222) & x(248) & x(249) & x(250) & x(276) & x(277) & x(278) & x(301) & x(302) & x(303) & x(305) & x(311) & x(326) & x(327) & x(328) & x(329) & x(330) & x(331) & x(353) & x(354) & x(356) & x(357) & x(358) & x(359) & x(400) & x(401) & x(412) & x(413) & x(414) & x(415) & x(416) & x(428) & x(429) & x(436) & x(441) & x(442) & x(443) & x(444) & x(450) & x(464) & x(469) & x(470) & x(471) & x(498) & x(507) & x(508) & x(514) & x(515) & x(523) & x(535) & x(536) & x(542) & x(543) & x(563) & x(564) & x(570) & x(571) & x(591) & x(597) & x(598) & x(619) & x(620) & x(647) & x(648) & x(649) & x(675) & x(676) & x(677) & x(678) & x(714) & x(715);
    y(205) <= not(p205_out);
    p205 : perceptron
        Generic map (
            WEIGHTS => "11111111110001000000000000011111111101111101111110011111111111111111111100",
            SHIFT => 4,
            B => 483,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p205_in,
            y(0) => p205_out,
            y(1 to 16 - 1) => dummy205
        );


    p206_in <= x(35) & x(37) & x(38) & x(39) & x(40) & x(41) & x(44) & x(45) & x(46) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(192) & x(194) & x(195) & x(220) & x(221) & x(222) & x(248) & x(249) & x(250) & x(276) & x(277) & x(278) & x(297) & x(298) & x(301) & x(302) & x(303) & x(305) & x(306) & x(325) & x(326) & x(327) & x(328) & x(329) & x(330) & x(331) & x(332) & x(346) & x(347) & x(348) & x(356) & x(357) & x(358) & x(359) & x(360) & x(373) & x(374) & x(375) & x(376) & x(400) & x(417) & x(438) & x(439) & x(450) & x(453) & x(466) & x(467) & x(479) & x(483) & x(484) & x(485) & x(487) & x(488) & x(494) & x(495) & x(496) & x(507) & x(513) & x(514) & x(515) & x(516) & x(518) & x(523) & x(535) & x(557) & x(563) & x(577) & x(605) & x(648) & x(649) & x(675) & x(676) & x(677) & x(678) & x(705) & x(709) & x(710) & x(766);
    y(206) <= not(p206_out);
    p206 : perceptron
        Generic map (
            WEIGHTS => "000000000000000000000000000000000111110011111111000111110000000001000111110000111110010000000000000",
            SHIFT => 4,
            B => -475,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p206_in,
            y(0) => p206_out,
            y(1 to 16 - 1) => dummy206
        );


    p207_in <= x(74) & x(75) & x(93) & x(94) & x(96) & x(103) & x(104) & x(105) & x(133) & x(166) & x(179) & x(182) & x(183) & x(207) & x(221) & x(239) & x(244) & x(248) & x(249) & x(250) & x(272) & x(274) & x(276) & x(277) & x(278) & x(303) & x(304) & x(305) & x(306) & x(334) & x(361) & x(362) & x(370) & x(371) & x(386) & x(387) & x(390) & x(398) & x(401) & x(413) & x(414) & x(418) & x(429) & x(445) & x(446) & x(473) & x(474) & x(500) & x(501) & x(502) & x(509) & x(528) & x(529) & x(556) & x(557) & x(558) & x(567) & x(568) & x(583) & x(584) & x(595) & x(607) & x(610) & x(611) & x(612) & x(627) & x(638) & x(640) & x(655) & x(656) & x(657) & x(685) & x(686) & x(717) & x(718) & x(720) & x(721) & x(748);
    y(207) <= not(p207_out);
    p207 : perceptron
        Generic map (
            WEIGHTS => "001110000111111111111111111111110000100001011111111111111111111111111111111111",
            SHIFT => 4,
            B => 729,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p207_in,
            y(0) => p207_out,
            y(1 to 16 - 1) => dummy207
        );


    p208_in <= x(37) & x(39) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(79) & x(93) & x(94) & x(95) & x(96) & x(102) & x(103) & x(104) & x(105) & x(106) & x(159) & x(192) & x(198) & x(199) & x(214) & x(226) & x(227) & x(239) & x(254) & x(265) & x(266) & x(267) & x(268) & x(270) & x(271) & x(272) & x(277) & x(283) & x(284) & x(294) & x(295) & x(296) & x(300) & x(303) & x(304) & x(309) & x(310) & x(311) & x(312) & x(320) & x(322) & x(323) & x(330) & x(338) & x(339) & x(361) & x(362) & x(366) & x(367) & x(373) & x(375) & x(376) & x(381) & x(382) & x(389) & x(390) & x(394) & x(403) & x(404) & x(409) & x(418) & x(431) & x(436) & x(458) & x(459) & x(460) & x(464) & x(488) & x(557) & x(659) & x(664) & x(665) & x(666) & x(667) & x(679) & x(693) & x(694) & x(695) & x(696) & x(708) & x(719) & x(720) & x(721) & x(722) & x(723) & x(736) & x(743) & x(748) & x(749) & x(764) & x(765) & x(769) & x(770) & x(771) & x(773) & x(774);
    y(208) <= not(p208_out);
    p208 : perceptron
        Generic map (
            WEIGHTS => "000000000000000000000000000010111111111111110111111111111011111111100000111000100000000100001000010000011001111111",
            SHIFT => 4,
            B => -140,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p208_in,
            y(0) => p208_out,
            y(1 to 16 - 1) => dummy208
        );


    p209_in <= x(37) & x(40) & x(45) & x(63) & x(64) & x(105) & x(108) & x(118) & x(124) & x(127) & x(146) & x(150) & x(151) & x(154) & x(164) & x(165) & x(181) & x(182) & x(191) & x(192) & x(193) & x(210) & x(219) & x(220) & x(221) & x(238) & x(247) & x(248) & x(249) & x(260) & x(261) & x(266) & x(276) & x(277) & x(289) & x(294) & x(295) & x(309) & x(319) & x(320) & x(323) & x(327) & x(330) & x(331) & x(332) & x(333) & x(338) & x(339) & x(346) & x(347) & x(348) & x(350) & x(361) & x(362) & x(366) & x(371) & x(373) & x(375) & x(389) & x(390) & x(391) & x(397) & x(403) & x(414) & x(418) & x(431) & x(444) & x(445) & x(446) & x(473) & x(474) & x(475) & x(479) & x(501) & x(502) & x(507) & x(528) & x(529) & x(535) & x(557) & x(558) & x(563) & x(584) & x(591) & x(619) & x(620) & x(640) & x(648) & x(661) & x(717) & x(718) & x(719) & x(720) & x(721) & x(723) & x(737) & x(738) & x(739) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(748) & x(750) & x(764) & x(769) & x(770) & x(773);
    y(209) <= not(p209_out);
    p209 : perceptron
        Generic map (
            WEIGHTS => "111111000000001100111011101111101110001100000000111000011100011101100000000000000000000010000000000000000000000",
            SHIFT => 4,
            B => -600,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p209_in,
            y(0) => p209_out,
            y(1 to 16 - 1) => dummy209
        );


    p210_in <= x(34) & x(35) & x(36) & x(37) & x(38) & x(39) & x(40) & x(41) & x(42) & x(44) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(79) & x(90) & x(91) & x(92) & x(93) & x(94) & x(95) & x(96) & x(97) & x(98) & x(99) & x(103) & x(104) & x(105) & x(106) & x(108) & x(135) & x(136) & x(155) & x(156) & x(163) & x(172) & x(192) & x(195) & x(242) & x(277) & x(292) & x(295) & x(304) & x(305) & x(323) & x(324) & x(333) & x(358) & x(359) & x(409) & x(418) & x(431) & x(437) & x(444) & x(446) & x(450) & x(458) & x(475) & x(485) & x(487) & x(507) & x(513) & x(514) & x(515) & x(516) & x(535) & x(541) & x(542) & x(543) & x(544) & x(563) & x(575) & x(584) & x(591) & x(612) & x(618) & x(619) & x(620) & x(647) & x(648) & x(675) & x(676) & x(677) & x(706) & x(707) & x(708) & x(709) & x(735) & x(737) & x(770) & x(777);
    y(210) <= not(p210_out);
    p210 : perceptron
        Generic map (
            WEIGHTS => "00000000000000000000000000000000000000000001100111111010111100110101101001000010000100101111111111111110",
            SHIFT => 4,
            B => -314,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p210_in,
            y(0) => p210_out,
            y(1 to 16 - 1) => dummy210
        );


    p211_in <= x(12) & x(37) & x(63) & x(64) & x(118) & x(124) & x(146) & x(192) & x(220) & x(248) & x(249) & x(291) & x(295) & x(296) & x(305) & x(306) & x(317) & x(320) & x(322) & x(323) & x(333) & x(342) & x(346) & x(347) & x(390) & x(418) & x(446) & x(450) & x(451) & x(473) & x(474) & x(475) & x(478) & x(479) & x(501) & x(502) & x(507) & x(529) & x(534) & x(535) & x(557) & x(558) & x(562) & x(563) & x(584) & x(591) & x(612) & x(618) & x(619) & x(620) & x(647) & x(648) & x(676) & x(731) & x(737) & x(738) & x(740) & x(741) & x(749) & x(750);
    y(211) <= not(p211_out);
    p211 : perceptron
        Generic map (
            WEIGHTS => "111100011111000011000111000000000000000000000000000001000000",
            SHIFT => 5,
            B => -832,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p211_in,
            y(0) => p211_out,
            y(1 to 17 - 1) => dummy211
        );


    p212_in <= x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(76) & x(77) & x(78) & x(79) & x(94) & x(95) & x(96) & x(103) & x(104) & x(105) & x(106) & x(107) & x(108) & x(192) & x(199) & x(221) & x(222) & x(227) & x(248) & x(249) & x(250) & x(277) & x(291) & x(301) & x(302) & x(303) & x(304) & x(318) & x(327) & x(328) & x(329) & x(330) & x(331) & x(332) & x(356) & x(357) & x(358) & x(359) & x(360) & x(433) & x(460) & x(473) & x(474) & x(485) & x(487) & x(488) & x(502) & x(513) & x(514) & x(515) & x(516) & x(542) & x(675) & x(676) & x(677) & x(678) & x(706) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(745) & x(746) & x(747) & x(748) & x(749) & x(764);
    y(212) <= not(p212_out);
    p212 : perceptron
        Generic map (
            WEIGHTS => "111111111111111111111000000000111111111111111111111111111111000001111111111110",
            SHIFT => 4,
            B => 602,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p212_in,
            y(0) => p212_out,
            y(1 to 16 - 1) => dummy212
        );


    p213_in <= x(98) & x(100) & x(108) & x(122) & x(124) & x(125) & x(152) & x(153) & x(163) & x(164) & x(165) & x(182) & x(183) & x(190) & x(191) & x(192) & x(193) & x(197) & x(210) & x(211) & x(220) & x(221) & x(222) & x(238) & x(248) & x(249) & x(277) & x(303) & x(304) & x(327) & x(328) & x(329) & x(330) & x(331) & x(332) & x(350) & x(356) & x(357) & x(358) & x(359) & x(463) & x(514) & x(515) & x(692) & x(693) & x(694) & x(695) & x(712) & x(715) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(724) & x(739) & x(740) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(748) & x(749);
    y(213) <= not(p213_out);
    p213 : perceptron
        Generic map (
            WEIGHTS => "111111110001100000110001000111111111111101111111111111111111111111111",
            SHIFT => 4,
            B => 462,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p213_in,
            y(0) => p213_out,
            y(1 to 16 - 1) => dummy213
        );


    p214_in <= x(69) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(104) & x(105) & x(135) & x(136) & x(163) & x(164) & x(165) & x(166) & x(192) & x(193) & x(194) & x(197) & x(220) & x(221) & x(222) & x(226) & x(238) & x(248) & x(249) & x(250) & x(266) & x(267) & x(276) & x(277) & x(278) & x(295) & x(300) & x(301) & x(302) & x(303) & x(305) & x(306) & x(320) & x(321) & x(329) & x(330) & x(331) & x(333) & x(334) & x(338) & x(346) & x(347) & x(348) & x(349) & x(350) & x(351) & x(358) & x(359) & x(360) & x(366) & x(375) & x(376) & x(377) & x(378) & x(450) & x(473) & x(474) & x(479) & x(481) & x(501) & x(502) & x(506) & x(507) & x(529) & x(534) & x(535) & x(556) & x(557) & x(558) & x(563) & x(584) & x(591) & x(611) & x(612) & x(638) & x(647) & x(648) & x(675) & x(676) & x(677) & x(679) & x(708) & x(719) & x(742) & x(743);
    y(214) <= not(p214_out);
    p214 : perceptron
        Generic map (
            WEIGHTS => "00000000000000000000001100011000111110000111001000000111100000110111001001110101110000000111",
            SHIFT => 4,
            B => -397,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p214_in,
            y(0) => p214_out,
            y(1 to 16 - 1) => dummy214
        );


    p215_in <= x(67) & x(68) & x(70) & x(109) & x(183) & x(198) & x(226) & x(227) & x(248) & x(249) & x(250) & x(254) & x(269) & x(275) & x(276) & x(277) & x(294) & x(295) & x(296) & x(297) & x(298) & x(303) & x(304) & x(306) & x(307) & x(309) & x(310) & x(311) & x(312) & x(320) & x(323) & x(324) & x(325) & x(331) & x(332) & x(334) & x(338) & x(339) & x(347) & x(348) & x(349) & x(352) & x(359) & x(360) & x(362) & x(366) & x(375) & x(376) & x(390) & x(394) & x(410) & x(414) & x(437) & x(442) & x(450) & x(461) & x(485) & x(486) & x(513) & x(514) & x(541) & x(542) & x(543) & x(656) & x(695) & x(696) & x(707) & x(709) & x(710) & x(711) & x(712) & x(720) & x(721) & x(722) & x(723) & x(735) & x(736) & x(737) & x(739) & x(741) & x(742) & x(743) & x(748) & x(749) & x(764) & x(765) & x(769) & x(770) & x(771) & x(772) & x(773) & x(774);
    y(215) <= not(p215_out);
    p215 : perceptron
        Generic map (
            WEIGHTS => "11101000111001110000011110000100011100111011101110010111111111111100000111100000001100000000",
            SHIFT => 4,
            B => 34,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p215_in,
            y(0) => p215_out,
            y(1 to 16 - 1) => dummy215
        );


    p216_in <= x(39) & x(40) & x(41) & x(43) & x(63) & x(66) & x(68) & x(69) & x(71) & x(105) & x(106) & x(107) & x(108) & x(151) & x(178) & x(179) & x(180) & x(184) & x(198) & x(209) & x(212) & x(220) & x(221) & x(226) & x(243) & x(248) & x(249) & x(250) & x(276) & x(277) & x(309) & x(310) & x(311) & x(324) & x(325) & x(326) & x(329) & x(338) & x(339) & x(346) & x(349) & x(355) & x(366) & x(375) & x(381) & x(383) & x(387) & x(388) & x(394) & x(416) & x(418) & x(437) & x(443) & x(444) & x(446) & x(450) & x(461) & x(462) & x(464) & x(473) & x(474) & x(475) & x(489) & x(490) & x(501) & x(502) & x(506) & x(518) & x(529) & x(530) & x(531) & x(537) & x(557) & x(564) & x(568) & x(569) & x(584) & x(592) & x(622) & x(625) & x(653) & x(654) & x(655) & x(675) & x(676) & x(677) & x(678) & x(703) & x(706) & x(707) & x(708) & x(709) & x(710) & x(714) & x(715) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(735) & x(736) & x(737) & x(738) & x(739) & x(740) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(764) & x(765) & x(769) & x(770) & x(771) & x(772) & x(773) & x(774);
    y(216) <= not(p216_out);
    p216 : perceptron
        Generic map (
            WEIGHTS => "11111111100001111101111011111100000000011001001101001101000000000010000101110111111111110000000000000000000000000000000000",
            SHIFT => 4,
            B => -328,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p216_in,
            y(0) => p216_out,
            y(1 to 17 - 1) => dummy216
        );


    p217_in <= x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(101) & x(102) & x(103) & x(104) & x(105) & x(106) & x(201) & x(256) & x(284) & x(291) & x(304) & x(309) & x(310) & x(311) & x(321) & x(322) & x(323) & x(331) & x(333) & x(338) & x(339) & x(342) & x(349) & x(350) & x(351) & x(361) & x(362) & x(366) & x(367) & x(369) & x(370) & x(371) & x(389) & x(390) & x(397) & x(398) & x(406) & x(417) & x(423) & x(425) & x(428) & x(433) & x(434) & x(445) & x(446) & x(451) & x(479) & x(507) & x(534) & x(535) & x(556) & x(562) & x(563) & x(591) & x(619) & x(647) & x(693) & x(694) & x(719) & x(721) & x(736) & x(748) & x(769);
    y(217) <= not(p217_out);
    p217 : perceptron
        Generic map (
            WEIGHTS => "111111111111111111011111111111011111110001100111001111111110111110000101",
            SHIFT => 4,
            B => 760,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p217_in,
            y(0) => p217_out,
            y(1 to 16 - 1) => dummy217
        );


    p218_in <= x(66) & x(67) & x(68) & x(73) & x(74) & x(94) & x(95) & x(97) & x(98) & x(105) & x(106) & x(107) & x(108) & x(129) & x(145) & x(156) & x(171) & x(172) & x(173) & x(180) & x(197) & x(199) & x(200) & x(201) & x(202) & x(227) & x(228) & x(242) & x(248) & x(249) & x(250) & x(255) & x(256) & x(276) & x(291) & x(294) & x(295) & x(296) & x(297) & x(299) & x(309) & x(311) & x(312) & x(322) & x(323) & x(324) & x(333) & x(339) & x(348) & x(351) & x(366) & x(390) & x(403) & x(409) & x(418) & x(422) & x(423) & x(431) & x(446) & x(450) & x(451) & x(458) & x(459) & x(474) & x(478) & x(479) & x(485) & x(486) & x(500) & x(501) & x(502) & x(506) & x(507) & x(514) & x(515) & x(526) & x(528) & x(529) & x(534) & x(535) & x(539) & x(542) & x(543) & x(544) & x(547) & x(548) & x(549) & x(553) & x(555) & x(557) & x(562) & x(563) & x(567) & x(568) & x(572) & x(579) & x(582) & x(584) & x(591) & x(610) & x(611) & x(612) & x(618) & x(619) & x(638) & x(647) & x(648) & x(649) & x(665) & x(666) & x(675) & x(676) & x(677) & x(678) & x(679) & x(680) & x(705) & x(706) & x(707) & x(708) & x(709) & x(732) & x(735) & x(736) & x(737) & x(743) & x(764) & x(765) & x(769) & x(770) & x(772) & x(773) & x(774);
    y(218) <= not(p218_out);
    p218 : perceptron
        Generic map (
            WEIGHTS => "0001100001111010111011111111000110011111111111110110010110011000110000011000001100000000001100000010001101110011111111111011111111111",
            SHIFT => 4,
            B => 339,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p218_in,
            y(0) => p218_out,
            y(1 to 17 - 1) => dummy218
        );


    p219_in <= x(62) & x(63) & x(64) & x(66) & x(68) & x(77) & x(78) & x(79) & x(104) & x(105) & x(106) & x(198) & x(199) & x(226) & x(227) & x(250) & x(254) & x(255) & x(256) & x(266) & x(267) & x(268) & x(282) & x(283) & x(284) & x(294) & x(295) & x(296) & x(309) & x(310) & x(311) & x(312) & x(322) & x(323) & x(338) & x(339) & x(347) & x(348) & x(349) & x(358) & x(359) & x(361) & x(362) & x(366) & x(367) & x(375) & x(376) & x(377) & x(386) & x(387) & x(388) & x(390) & x(403) & x(404) & x(405) & x(409) & x(414) & x(418) & x(424) & x(432) & x(433) & x(446) & x(460) & x(474) & x(487) & x(647) & x(690) & x(693) & x(694) & x(695) & x(719) & x(720) & x(721) & x(722) & x(723) & x(736) & x(742) & x(743) & x(744) & x(748) & x(764) & x(765) & x(766) & x(769) & x(770) & x(771) & x(772) & x(773) & x(774);
    y(219) <= not(p219_out);
    p219 : perceptron
        Generic map (
            WEIGHTS => "11111111111000000000000000000000000011111000011111101111101110101111111111100001000000000",
            SHIFT => 4,
            B => -139,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p219_in,
            y(0) => p219_out,
            y(1 to 16 - 1) => dummy219
        );


    p220_in <= x(40) & x(108) & x(163) & x(182) & x(183) & x(191) & x(192) & x(193) & x(210) & x(211) & x(212) & x(219) & x(220) & x(221) & x(237) & x(238) & x(239) & x(247) & x(248) & x(249) & x(266) & x(275) & x(277) & x(303) & x(320) & x(323) & x(328) & x(329) & x(330) & x(331) & x(332) & x(350) & x(358) & x(390) & x(416) & x(418) & x(446) & x(473) & x(474) & x(475) & x(501) & x(502) & x(514) & x(515) & x(529) & x(557) & x(704) & x(709) & x(711) & x(712) & x(713) & x(715) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(737) & x(738) & x(739) & x(740) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(748) & x(749);
    y(220) <= not(p220_out);
    p220 : perceptron
        Generic map (
            WEIGHTS => "0101100011100011100010010111111111011111111111011111111111111111111111111",
            SHIFT => 4,
            B => 566,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p220_in,
            y(0) => p220_out,
            y(1 to 16 - 1) => dummy220
        );


    p221_in <= x(34) & x(35) & x(36) & x(37) & x(38) & x(39) & x(40) & x(41) & x(45) & x(46) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(79) & x(101) & x(102) & x(103) & x(104) & x(105) & x(106) & x(107) & x(108) & x(118) & x(151) & x(187) & x(216) & x(218) & x(222) & x(249) & x(250) & x(268) & x(269) & x(277) & x(317) & x(327) & x(330) & x(343) & x(344) & x(348) & x(355) & x(357) & x(358) & x(362) & x(379) & x(380) & x(386) & x(387) & x(390) & x(394) & x(407) & x(414) & x(415) & x(418) & x(431) & x(432) & x(446) & x(453) & x(473) & x(474) & x(486) & x(487) & x(495) & x(500) & x(501) & x(502) & x(513) & x(514) & x(515) & x(528) & x(529) & x(530) & x(535) & x(536) & x(556) & x(557) & x(558) & x(564) & x(566) & x(579) & x(580) & x(583) & x(584) & x(585) & x(591) & x(597) & x(611) & x(612) & x(613) & x(620) & x(637) & x(638) & x(640) & x(648) & x(649) & x(691) & x(692) & x(693) & x(703) & x(720) & x(721) & x(722);
    y(221) <= not(p221_out);
    p221 : perceptron
        Generic map (
            WEIGHTS => "1111111111111111111111111111111111110000000000011111111101111011110110000110000111000000000000000000000000001110111",
            SHIFT => 4,
            B => 184,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p221_in,
            y(0) => p221_out,
            y(1 to 16 - 1) => dummy221
        );


    p222_in <= x(35) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(97) & x(101) & x(102) & x(103) & x(104) & x(105) & x(106) & x(107) & x(108) & x(122) & x(125) & x(162) & x(163) & x(164) & x(165) & x(171) & x(190) & x(191) & x(192) & x(193) & x(199) & x(200) & x(210) & x(211) & x(218) & x(219) & x(220) & x(221) & x(222) & x(246) & x(247) & x(248) & x(249) & x(250) & x(272) & x(273) & x(274) & x(276) & x(277) & x(294) & x(309) & x(323) & x(327) & x(329) & x(330) & x(331) & x(332) & x(338) & x(357) & x(358) & x(359) & x(417) & x(450) & x(506) & x(507) & x(528) & x(556) & x(584) & x(611) & x(638) & x(656) & x(659) & x(686) & x(695) & x(697) & x(706) & x(707) & x(708) & x(709) & x(710) & x(711) & x(712) & x(713) & x(714) & x(715) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(734) & x(735) & x(736) & x(737) & x(738) & x(739) & x(740) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(748) & x(749) & x(770) & x(772);
    y(222) <= not(p222_out);
    p222 : perceptron
        Generic map (
            WEIGHTS => "000000000000000000000000111101111000011111111111111100000000000000001111111101000000000000000000000000000000000000",
            SHIFT => 5,
            B => -1083,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p222_in,
            y(0) => p222_out,
            y(1 to 17 - 1) => dummy222
        );


    p223_in <= x(66) & x(67) & x(69) & x(138) & x(165) & x(166) & x(193) & x(194) & x(201) & x(202) & x(210) & x(211) & x(220) & x(221) & x(222) & x(231) & x(232) & x(248) & x(249) & x(250) & x(256) & x(257) & x(265) & x(276) & x(277) & x(278) & x(297) & x(299) & x(305) & x(306) & x(309) & x(310) & x(311) & x(333) & x(334) & x(337) & x(349) & x(350) & x(351) & x(360) & x(366) & x(376) & x(377) & x(378) & x(405) & x(406) & x(422) & x(433) & x(482) & x(511) & x(512) & x(529) & x(545) & x(555) & x(557) & x(584) & x(614) & x(670) & x(693) & x(694) & x(695) & x(704) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(724) & x(747) & x(748) & x(749);
    y(223) <= not(p223_out);
    p223 : perceptron
        Generic map (
            WEIGHTS => "0000000011000001100011100011001110010001100000101111111111000100000000000",
            SHIFT => 4,
            B => -311,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p223_in,
            y(0) => p223_out,
            y(1 to 16 - 1) => dummy223
        );


    p224_in <= x(37) & x(38) & x(39) & x(40) & x(41) & x(45) & x(46) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(79) & x(102) & x(103) & x(104) & x(105) & x(106) & x(135) & x(192) & x(198) & x(215) & x(249) & x(267) & x(277) & x(301) & x(302) & x(303) & x(304) & x(309) & x(329) & x(330) & x(331) & x(332) & x(338) & x(339) & x(347) & x(348) & x(361) & x(362) & x(366) & x(370) & x(371) & x(373) & x(375) & x(386) & x(387) & x(388) & x(389) & x(390) & x(396) & x(398) & x(399) & x(400) & x(401) & x(402) & x(413) & x(414) & x(415) & x(416) & x(418) & x(437) & x(446) & x(450) & x(473) & x(474) & x(475) & x(501) & x(502) & x(528) & x(529) & x(556) & x(557) & x(558) & x(582) & x(640) & x(641) & x(648) & x(675) & x(676) & x(677) & x(678) & x(705) & x(739) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747);
    y(224) <= not(p224_out);
    p224 : perceptron
        Generic map (
            WEIGHTS => "111111111111111111111111111111110010100000000000110001111111001111111111010100000000000001111110000000",
            SHIFT => 4,
            B => 341,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p224_in,
            y(0) => p224_out,
            y(1 to 16 - 1) => dummy224
        );


    p225_in <= x(40) & x(68) & x(100) & x(107) & x(108) & x(123) & x(145) & x(162) & x(172) & x(221) & x(222) & x(240) & x(241) & x(248) & x(249) & x(250) & x(268) & x(276) & x(277) & x(278) & x(295) & x(297) & x(298) & x(299) & x(302) & x(303) & x(323) & x(325) & x(326) & x(327) & x(328) & x(329) & x(330) & x(331) & x(350) & x(357) & x(400) & x(416) & x(430) & x(431) & x(457) & x(458) & x(459) & x(483) & x(498) & x(510) & x(540) & x(541) & x(542) & x(543) & x(544) & x(549) & x(550) & x(552) & x(568) & x(571) & x(572) & x(657) & x(716) & x(740) & x(742) & x(743) & x(744) & x(745);
    y(225) <= not(p225_out);
    p225 : perceptron
        Generic map (
            WEIGHTS => "1110010101100111011100000000000000001111111111111111111110000000",
            SHIFT => 4,
            B => 36,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p225_in,
            y(0) => p225_out,
            y(1 to 16 - 1) => dummy225
        );


    p226_in <= x(34) & x(35) & x(36) & x(37) & x(38) & x(39) & x(40) & x(41) & x(42) & x(43) & x(44) & x(45) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(79) & x(90) & x(91) & x(92) & x(93) & x(94) & x(95) & x(96) & x(97) & x(98) & x(99) & x(100) & x(101) & x(102) & x(103) & x(104) & x(105) & x(106) & x(107) & x(108) & x(163) & x(164) & x(191) & x(192) & x(193) & x(198) & x(226) & x(249) & x(254) & x(265) & x(266) & x(267) & x(277) & x(279) & x(292) & x(293) & x(294) & x(303) & x(305) & x(309) & x(310) & x(311) & x(329) & x(330) & x(331) & x(334) & x(337) & x(338) & x(339) & x(357) & x(358) & x(366) & x(367) & x(369) & x(371) & x(394) & x(396) & x(397) & x(398) & x(399) & x(400) & x(417) & x(424) & x(425) & x(428) & x(445) & x(450) & x(453) & x(487) & x(514) & x(515) & x(516) & x(534) & x(535) & x(542) & x(543) & x(544) & x(647) & x(675) & x(693) & x(694) & x(703) & x(707) & x(715) & x(716) & x(717) & x(718) & x(719) & x(720) & x(734) & x(735) & x(736) & x(737) & x(738) & x(739) & x(740) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(750) & x(761) & x(763) & x(764) & x(765) & x(766) & x(769) & x(770) & x(771) & x(772) & x(773) & x(774) & x(775);
    y(226) <= not(p226_out);
    p226 : perceptron
        Generic map (
            WEIGHTS => "1111111111111111111111111111111111111111111111111000001101111001111011111101111111001000001000100111100111000001111111111111111111111111111111111",
            SHIFT => 4,
            B => 1330,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p226_in,
            y(0) => p226_out,
            y(1 to 17 - 1) => dummy226
        );


    p227_in <= x(35) & x(37) & x(38) & x(39) & x(40) & x(41) & x(42) & x(43) & x(46) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(79) & x(91) & x(92) & x(94) & x(96) & x(97) & x(98) & x(99) & x(100) & x(102) & x(103) & x(104) & x(105) & x(106) & x(108) & x(163) & x(171) & x(172) & x(197) & x(211) & x(226) & x(248) & x(249) & x(250) & x(254) & x(276) & x(292) & x(295) & x(296) & x(297) & x(305) & x(311) & x(323) & x(324) & x(331) & x(359) & x(418) & x(422) & x(423) & x(425) & x(446) & x(450) & x(473) & x(474) & x(475) & x(487) & x(502) & x(507) & x(513) & x(514) & x(515) & x(516) & x(529) & x(530) & x(531) & x(534) & x(535) & x(541) & x(542) & x(543) & x(544) & x(557) & x(558) & x(563) & x(571) & x(591) & x(618) & x(619) & x(648) & x(676) & x(692) & x(695) & x(715) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(740) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(748) & x(749);
    y(227) <= not(p227_out);
    p227 : perceptron
        Generic map (
            WEIGHTS => "000000000000000000000000000000000000000001111000000001111111001111111110110000111110000111011111000000000000000000000",
            SHIFT => 4,
            B => -719,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p227_in,
            y(0) => p227_out,
            y(1 to 16 - 1) => dummy227
        );


    p228_in <= x(40) & x(67) & x(68) & x(69) & x(70) & x(105) & x(109) & x(138) & x(166) & x(193) & x(198) & x(211) & x(212) & x(248) & x(249) & x(250) & x(271) & x(276) & x(277) & x(278) & x(299) & x(304) & x(306) & x(309) & x(324) & x(325) & x(326) & x(327) & x(334) & x(352) & x(362) & x(380) & x(391) & x(394) & x(404) & x(409) & x(436) & x(437) & x(444) & x(464) & x(465) & x(540) & x(541) & x(542) & x(543) & x(544) & x(545) & x(571) & x(572) & x(573) & x(574) & x(706) & x(707) & x(708) & x(716) & x(735) & x(736) & x(737) & x(739) & x(742) & x(743) & x(744) & x(745) & x(746) & x(773);
    y(228) <= not(p228_out);
    p228 : perceptron
        Generic map (
            WEIGHTS => "11111001110001110111011000001010100000100111111111100000000000000",
            SHIFT => 4,
            B => 43,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p228_in,
            y(0) => p228_out,
            y(1 to 16 - 1) => dummy228
        );


    p229_in <= x(35) & x(37) & x(38) & x(39) & x(40) & x(41) & x(45) & x(46) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(78) & x(79) & x(102) & x(104) & x(105) & x(118) & x(192) & x(198) & x(208) & x(211) & x(221) & x(222) & x(249) & x(277) & x(302) & x(303) & x(309) & x(325) & x(326) & x(328) & x(329) & x(330) & x(331) & x(332) & x(338) & x(339) & x(350) & x(362) & x(366) & x(371) & x(387) & x(390) & x(394) & x(400) & x(402) & x(412) & x(414) & x(415) & x(416) & x(418) & x(446) & x(450) & x(473) & x(474) & x(475) & x(501) & x(502) & x(514) & x(528) & x(529) & x(530) & x(531) & x(557) & x(558) & x(584) & x(612) & x(640) & x(675) & x(676) & x(677) & x(678) & x(703) & x(707) & x(709) & x(714) & x(715) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(736) & x(737) & x(738) & x(739) & x(740) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(748) & x(749) & x(750) & x(764) & x(770) & x(771) & x(772) & x(773) & x(774) & x(775);
    y(229) <= not(p229_out);
    p229 : perceptron
        Generic map (
            WEIGHTS => "00000000000000000000000000001011100001111111111110110011000000110111111111111111000001111111111111111111111111111111111",
            SHIFT => 5,
            B => 528,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p229_in,
            y(0) => p229_out,
            y(1 to 18 - 1) => dummy229
        );


    p230_in <= x(125) & x(126) & x(153) & x(154) & x(161) & x(171) & x(172) & x(191) & x(192) & x(200) & x(228) & x(248) & x(264) & x(266) & x(267) & x(288) & x(289) & x(290) & x(292) & x(304) & x(317) & x(318) & x(322) & x(323) & x(330) & x(331) & x(332) & x(333) & x(343) & x(344) & x(348) & x(350) & x(361) & x(362) & x(368) & x(378) & x(389) & x(404) & x(433) & x(450) & x(478) & x(479) & x(507) & x(524) & x(534) & x(535) & x(537) & x(552) & x(553) & x(563) & x(565) & x(591) & x(593) & x(619) & x(646) & x(647) & x(648);
    y(230) <= not(p230_out);
    p230 : perceptron
        Generic map (
            WEIGHTS => "000010011001100111101100000011100010010000000000000000000",
            SHIFT => 4,
            B => -422,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p230_in,
            y(0) => p230_out,
            y(1 to 15 - 1) => dummy230
        );


    p231_in <= x(3) & x(4) & x(7) & x(8) & x(10) & x(19) & x(23) & x(24) & x(28) & x(35) & x(53) & x(54) & x(57) & x(58) & x(61) & x(75) & x(76) & x(79) & x(84) & x(104) & x(108) & x(110) & x(124) & x(125) & x(142) & x(151) & x(153) & x(155) & x(163) & x(164) & x(165) & x(166) & x(171) & x(172) & x(173) & x(181) & x(182) & x(191) & x(192) & x(193) & x(194) & x(196) & x(197) & x(198) & x(199) & x(200) & x(201) & x(214) & x(215) & x(219) & x(220) & x(221) & x(226) & x(227) & x(228) & x(239) & x(248) & x(249) & x(250) & x(254) & x(255) & x(256) & x(266) & x(267) & x(268) & x(276) & x(277) & x(283) & x(288) & x(290) & x(294) & x(295) & x(296) & x(297) & x(298) & x(309) & x(310) & x(311) & x(315) & x(316) & x(317) & x(320) & x(322) & x(323) & x(332) & x(334) & x(338) & x(339) & x(346) & x(347) & x(348) & x(349) & x(364) & x(366) & x(375) & x(376) & x(380) & x(381) & x(392) & x(403) & x(408) & x(419) & x(431) & x(433) & x(436) & x(448) & x(450) & x(459) & x(460) & x(474) & x(479) & x(501) & x(502) & x(503) & x(507) & x(509) & x(529) & x(534) & x(535) & x(537) & x(557) & x(562) & x(563) & x(564) & x(565) & x(584) & x(591) & x(592) & x(612) & x(619) & x(620) & x(622) & x(624) & x(625) & x(643) & x(644) & x(647) & x(648) & x(662) & x(664) & x(671) & x(673) & x(675) & x(676) & x(677) & x(678) & x(679) & x(692) & x(693) & x(705) & x(706) & x(707) & x(708) & x(709) & x(710) & x(711) & x(712) & x(725) & x(729) & x(735) & x(736) & x(737) & x(738) & x(739) & x(740) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(750) & x(760) & x(763) & x(764) & x(765) & x(766) & x(768) & x(769) & x(770) & x(771) & x(772) & x(773) & x(774) & x(775) & x(779);
    y(231) <= not(p231_out);
    p231 : perceptron
        Generic map (
            WEIGHTS => "1111111110111111101101001000111100000111110000000111000011100000011011000000001111000100111110111111111111011000010000000000000000000011001111000001100000000110000000000000010000000000001",
            SHIFT => 4,
            B => 484,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p231_in,
            y(0) => p231_out,
            y(1 to 17 - 1) => dummy231
        );


    p232_in <= x(39) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(77) & x(91) & x(92) & x(93) & x(94) & x(104) & x(105) & x(152) & x(153) & x(171) & x(179) & x(180) & x(181) & x(193) & x(247) & x(248) & x(249) & x(254) & x(276) & x(277) & x(291) & x(292) & x(295) & x(322) & x(323) & x(324) & x(350) & x(351) & x(367) & x(378) & x(450) & x(507) & x(535) & x(563) & x(624) & x(625) & x(675) & x(677);
    y(232) <= not(p232_out);
    p232 : perceptron
        Generic map (
            WEIGHTS => "000000000000000001111110000000001111110111111111",
            SHIFT => 4,
            B => -294,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p232_in,
            y(0) => p232_out,
            y(1 to 15 - 1) => dummy232
        );


    p233_in <= x(35) & x(37) & x(39) & x(40) & x(44) & x(62) & x(63) & x(64) & x(66) & x(67) & x(68) & x(69) & x(70) & x(72) & x(77) & x(78) & x(79) & x(90) & x(104) & x(105) & x(106) & x(107) & x(108) & x(136) & x(163) & x(164) & x(184) & x(185) & x(186) & x(230) & x(231) & x(232) & x(257) & x(258) & x(259) & x(260) & x(284) & x(298) & x(321) & x(326) & x(330) & x(331) & x(338) & x(353) & x(354) & x(358) & x(360) & x(367) & x(369) & x(370) & x(378) & x(396) & x(397) & x(398) & x(400) & x(401) & x(402) & x(414) & x(416) & x(425) & x(427) & x(428) & x(429) & x(430) & x(436) & x(437) & x(444) & x(446) & x(456) & x(457) & x(491) & x(501) & x(502) & x(515) & x(516) & x(528) & x(529) & x(530) & x(542) & x(543) & x(544) & x(556) & x(557) & x(569) & x(584) & x(612);
    y(233) <= not(p233_out);
    p233 : perceptron
        Generic map (
            WEIGHTS => "11111111111111111111111000000111111111111111110100000000000000001100001001100011100000",
            SHIFT => 4,
            B => 181,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p233_in,
            y(0) => p233_out,
            y(1 to 16 - 1) => dummy233
        );


    p234_in <= x(35) & x(39) & x(40) & x(41) & x(44) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(79) & x(90) & x(91) & x(92) & x(93) & x(94) & x(95) & x(96) & x(97) & x(98) & x(100) & x(102) & x(105) & x(106) & x(108) & x(136) & x(145) & x(191) & x(192) & x(193) & x(209) & x(211) & x(212) & x(213) & x(220) & x(235) & x(236) & x(237) & x(238) & x(239) & x(240) & x(241) & x(242) & x(263) & x(266) & x(270) & x(271) & x(272) & x(273) & x(299) & x(300) & x(305) & x(323) & x(328) & x(333) & x(334) & x(338) & x(349) & x(350) & x(359) & x(361) & x(366) & x(376) & x(377) & x(378) & x(388) & x(406) & x(423) & x(433) & x(434) & x(445) & x(450) & x(461) & x(462) & x(473) & x(489) & x(490) & x(501) & x(514) & x(517) & x(529) & x(535) & x(542) & x(543) & x(545) & x(557) & x(627) & x(628) & x(638) & x(656) & x(657) & x(693) & x(732) & x(738) & x(739) & x(740) & x(741) & x(742) & x(743);
    y(234) <= not(p234_out);
    p234 : perceptron
        Generic map (
            WEIGHTS => "00000000000000000000000000000011111000010000000000000000110110110101110111101110110010100100000010000000",
            SHIFT => 3,
            B => -379,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p234_in,
            y(0) => p234_out,
            y(1 to 15 - 1) => dummy234
        );


    p235_in <= x(34) & x(35) & x(36) & x(37) & x(38) & x(39) & x(40) & x(41) & x(45) & x(46) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(79) & x(102) & x(103) & x(104) & x(105) & x(106) & x(107) & x(108) & x(118) & x(123) & x(124) & x(125) & x(146) & x(147) & x(152) & x(154) & x(155) & x(163) & x(174) & x(184) & x(185) & x(190) & x(191) & x(210) & x(260) & x(295) & x(302) & x(303) & x(305) & x(317) & x(323) & x(330) & x(331) & x(333) & x(338) & x(339) & x(342) & x(347) & x(348) & x(361) & x(362) & x(371) & x(373) & x(375) & x(378) & x(386) & x(387) & x(388) & x(390) & x(398) & x(406) & x(414) & x(415) & x(416) & x(418) & x(433) & x(440) & x(441) & x(444) & x(446) & x(460) & x(473) & x(474) & x(475) & x(479) & x(500) & x(501) & x(502) & x(507) & x(528) & x(529) & x(530) & x(535) & x(537) & x(555) & x(556) & x(557) & x(558) & x(563) & x(565) & x(566) & x(567) & x(583) & x(584) & x(585) & x(591) & x(594) & x(602) & x(611) & x(612) & x(613) & x(619) & x(638) & x(639) & x(640) & x(695) & x(719) & x(721) & x(722) & x(769);
    y(235) <= not(p235_out);
    p235 : perceptron
        Generic map (
            WEIGHTS => "1111111111111111111111111111111111100000000010001101000010000001110011101110101110011100000000000000000000000000001000000011110",
            SHIFT => 4,
            B => 14,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p235_in,
            y(0) => p235_out,
            y(1 to 17 - 1) => dummy235
        );


    p236_in <= x(35) & x(43) & x(66) & x(68) & x(69) & x(73) & x(165) & x(166) & x(192) & x(193) & x(194) & x(220) & x(221) & x(248) & x(249) & x(250) & x(276) & x(277) & x(278) & x(297) & x(302) & x(305) & x(306) & x(309) & x(310) & x(311) & x(321) & x(322) & x(326) & x(329) & x(330) & x(333) & x(334) & x(337) & x(338) & x(348) & x(349) & x(350) & x(351) & x(357) & x(358) & x(361) & x(362) & x(366) & x(376) & x(377) & x(378) & x(379) & x(394) & x(405) & x(406) & x(425) & x(433) & x(450) & x(454) & x(455) & x(473) & x(474) & x(501) & x(502) & x(506) & x(507) & x(528) & x(529) & x(530) & x(556) & x(557) & x(584) & x(612) & x(647) & x(674) & x(720) & x(742) & x(743) & x(744) & x(769) & x(770) & x(773);
    y(236) <= not(p236_out);
    p236 : perceptron
        Generic map (
            WEIGHTS => "111111111111111111100110001100011001111001101111011011000000110000000111000000",
            SHIFT => 4,
            B => 54,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p236_in,
            y(0) => p236_out,
            y(1 to 16 - 1) => dummy236
        );


    p237_in <= x(35) & x(38) & x(39) & x(40) & x(41) & x(43) & x(44) & x(49) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(79) & x(90) & x(91) & x(92) & x(93) & x(94) & x(95) & x(96) & x(97) & x(98) & x(99) & x(102) & x(103) & x(104) & x(105) & x(106) & x(210) & x(221) & x(222) & x(248) & x(249) & x(250) & x(276) & x(277) & x(278) & x(296) & x(297) & x(298) & x(299) & x(300) & x(301) & x(302) & x(303) & x(305) & x(306) & x(325) & x(326) & x(329) & x(330) & x(331) & x(332) & x(357) & x(358) & x(359) & x(360) & x(417) & x(425) & x(446) & x(450) & x(453) & x(454) & x(479) & x(483) & x(507) & x(513) & x(530) & x(535) & x(557) & x(558) & x(647) & x(648) & x(649) & x(675) & x(676) & x(677) & x(695) & x(711) & x(712) & x(717) & x(718) & x(719) & x(720) & x(721) & x(723) & x(747) & x(748);
    y(237) <= not(p237_out);
    p237 : perceptron
        Generic map (
            WEIGHTS => "11111111111111111111111111111111111111111111111111000000001100000000001001001010010011111111111111111",
            SHIFT => 4,
            B => 1114,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p237_in,
            y(0) => p237_out,
            y(1 to 16 - 1) => dummy237
        );


    p238_in <= x(37) & x(63) & x(64) & x(65) & x(66) & x(68) & x(70) & x(74) & x(78) & x(79) & x(95) & x(98) & x(99) & x(100) & x(101) & x(102) & x(103) & x(104) & x(105) & x(106) & x(181) & x(182) & x(190) & x(210) & x(211) & x(212) & x(231) & x(255) & x(257) & x(259) & x(275) & x(284) & x(307) & x(361) & x(362) & x(390) & x(416) & x(418) & x(434) & x(444) & x(446) & x(450) & x(463) & x(490) & x(491) & x(507) & x(515) & x(518) & x(535) & x(563) & x(591) & x(592) & x(619) & x(620) & x(622) & x(647) & x(648) & x(675) & x(676) & x(677) & x(693) & x(694) & x(709) & x(712) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(723) & x(732) & x(746) & x(747) & x(748) & x(749);
    y(238) <= not(p238_out);
    p238 : perceptron
        Generic map (
            WEIGHTS => "1111111111111111111111011100000000001001010001001111111111111111111111111111",
            SHIFT => 5,
            B => 893,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p238_in,
            y(0) => p238_out,
            y(1 to 17 - 1) => dummy238
        );


    p239_in <= x(35) & x(37) & x(38) & x(39) & x(40) & x(41) & x(45) & x(46) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(78) & x(79) & x(102) & x(103) & x(104) & x(105) & x(108) & x(164) & x(192) & x(198) & x(211) & x(212) & x(221) & x(222) & x(226) & x(236) & x(237) & x(239) & x(240) & x(249) & x(261) & x(263) & x(264) & x(277) & x(298) & x(299) & x(300) & x(301) & x(302) & x(303) & x(304) & x(309) & x(311) & x(326) & x(327) & x(328) & x(329) & x(330) & x(331) & x(332) & x(337) & x(338) & x(339) & x(350) & x(357) & x(358) & x(361) & x(362) & x(366) & x(378) & x(390) & x(394) & x(398) & x(400) & x(401) & x(406) & x(411) & x(414) & x(416) & x(418) & x(434) & x(438) & x(446) & x(450) & x(461) & x(462) & x(473) & x(474) & x(475) & x(486) & x(489) & x(501) & x(502) & x(506) & x(507) & x(514) & x(528) & x(529) & x(531) & x(535) & x(544) & x(557) & x(558) & x(573) & x(640) & x(647) & x(648) & x(649) & x(675) & x(676) & x(677) & x(678) & x(687) & x(703) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(736) & x(737) & x(738) & x(739) & x(740) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(770) & x(773);
    y(239) <= not(p239_out);
    p239 : perceptron
        Generic map (
            WEIGHTS => "1111111111111111111111111111011000110000010001000000000000000000010000010011111110110111000110011000011001011111110100000000000000000000",
            SHIFT => 4,
            B => -64,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p239_in,
            y(0) => p239_out,
            y(1 to 17 - 1) => dummy239
        );


    p240_in <= x(35) & x(37) & x(39) & x(40) & x(41) & x(43) & x(46) & x(47) & x(63) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(77) & x(78) & x(107) & x(108) & x(163) & x(191) & x(192) & x(193) & x(199) & x(207) & x(221) & x(227) & x(248) & x(249) & x(266) & x(277) & x(293) & x(294) & x(295) & x(305) & x(306) & x(309) & x(322) & x(331) & x(334) & x(338) & x(348) & x(359) & x(360) & x(366) & x(376) & x(386) & x(387) & x(388) & x(414) & x(415) & x(416) & x(432) & x(433) & x(444) & x(446) & x(456) & x(460) & x(464) & x(473) & x(474) & x(475) & x(488) & x(501) & x(502) & x(528) & x(529) & x(530) & x(531) & x(543) & x(544) & x(556) & x(557) & x(558) & x(566) & x(567) & x(568) & x(583) & x(584) & x(594) & x(595) & x(606) & x(611) & x(612) & x(634) & x(636) & x(637) & x(638) & x(640) & x(656) & x(666) & x(667) & x(677) & x(706) & x(741) & x(742) & x(743) & x(746) & x(747);
    y(240) <= not(p240_out);
    p240 : perceptron
        Generic map (
            WEIGHTS => "1111111111111111111111100001001001011100111010111011111100101000000000000110000000000000000000001111111",
            SHIFT => 4,
            B => 119,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p240_in,
            y(0) => p240_out,
            y(1 to 16 - 1) => dummy240
        );


    p241_in <= x(35) & x(37) & x(38) & x(39) & x(40) & x(41) & x(42) & x(43) & x(45) & x(46) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(79) & x(98) & x(99) & x(100) & x(101) & x(102) & x(103) & x(104) & x(105) & x(106) & x(107) & x(108) & x(150) & x(155) & x(178) & x(179) & x(210) & x(218) & x(221) & x(248) & x(249) & x(250) & x(276) & x(277) & x(305) & x(306) & x(347) & x(348) & x(362) & x(376) & x(418) & x(446) & x(450) & x(453) & x(474) & x(478) & x(479) & x(481) & x(490) & x(494) & x(501) & x(502) & x(506) & x(507) & x(517) & x(528) & x(529) & x(530) & x(534) & x(535) & x(556) & x(557) & x(558) & x(563) & x(583) & x(584) & x(586) & x(591) & x(611) & x(612) & x(619) & x(638) & x(647) & x(648) & x(649) & x(675) & x(676) & x(677) & x(678) & x(679) & x(680) & x(681) & x(693) & x(694) & x(695) & x(705) & x(706) & x(707) & x(708) & x(709) & x(710) & x(711) & x(712) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(724) & x(733) & x(734) & x(736) & x(737) & x(739) & x(740) & x(742) & x(744) & x(745) & x(746) & x(747) & x(748) & x(749);
    y(241) <= not(p241_out);
    p241 : perceptron
        Generic map (
            WEIGHTS => "111111111111111111111111111111111111111101110111111111101001001100100110000110001000100101111111111111111111111111111111111111111111",
            SHIFT => 5,
            B => 2111,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p241_in,
            y(0) => p241_out,
            y(1 to 18 - 1) => dummy241
        );


    p242_in <= x(38) & x(39) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(72) & x(73) & x(74) & x(75) & x(78) & x(79) & x(102) & x(103) & x(104) & x(105) & x(106) & x(118) & x(151) & x(152) & x(155) & x(172) & x(173) & x(174) & x(182) & x(200) & x(202) & x(270) & x(277) & x(295) & x(317) & x(320) & x(327) & x(332) & x(333) & x(342) & x(343) & x(361) & x(362) & x(390) & x(418) & x(446) & x(450) & x(458) & x(474) & x(475) & x(479) & x(502) & x(507) & x(509) & x(525) & x(534) & x(535) & x(551) & x(557) & x(562) & x(563) & x(564) & x(565) & x(566) & x(580) & x(591) & x(593) & x(594) & x(619) & x(622) & x(625) & x(640) & x(647) & x(719) & x(721) & x(738) & x(769);
    y(242) <= not(p242_out);
    p242 : perceptron
        Generic map (
            WEIGHTS => "111111111111111111111100000000000101100011000000100000000000000000000000001100",
            SHIFT => 5,
            B => -285,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p242_in,
            y(0) => p242_out,
            y(1 to 17 - 1) => dummy242
        );


    p243_in <= x(138) & x(166) & x(193) & x(198) & x(217) & x(221) & x(226) & x(244) & x(247) & x(248) & x(249) & x(250) & x(275) & x(276) & x(277) & x(278) & x(294) & x(295) & x(304) & x(305) & x(306) & x(307) & x(309) & x(310) & x(311) & x(320) & x(332) & x(333) & x(334) & x(338) & x(339) & x(346) & x(347) & x(348) & x(349) & x(361) & x(366) & x(375) & x(376) & x(378) & x(386) & x(387) & x(394) & x(414) & x(415) & x(443) & x(450) & x(469) & x(489) & x(495) & x(506) & x(517) & x(518) & x(534) & x(535) & x(562) & x(591) & x(619) & x(627) & x(646) & x(647) & x(648) & x(655) & x(656) & x(657) & x(658) & x(660) & x(674) & x(675) & x(695) & x(712) & x(736) & x(737) & x(739) & x(740) & x(741) & x(742) & x(743) & x(744) & x(764) & x(765) & x(769) & x(770) & x(772) & x(773);
    y(243) <= not(p243_out);
    p243 : perceptron
        Generic map (
            WEIGHTS => "1110110111111111001111000111100111110110110111110110011111111111111111000000000000000",
            SHIFT => 4,
            B => 295,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p243_in,
            y(0) => p243_out,
            y(1 to 16 - 1) => dummy243
        );


    p244_in <= x(0) & x(1) & x(2) & x(3) & x(4) & x(5) & x(6) & x(7) & x(8) & x(9) & x(10) & x(11) & x(12) & x(15) & x(16) & x(17) & x(18) & x(19) & x(20) & x(21) & x(22) & x(23) & x(24) & x(25) & x(26) & x(27) & x(28) & x(29) & x(30) & x(31) & x(32) & x(33) & x(34) & x(35) & x(36) & x(37) & x(38) & x(39) & x(40) & x(41) & x(42) & x(43) & x(44) & x(45) & x(46) & x(52) & x(53) & x(54) & x(55) & x(56) & x(57) & x(58) & x(59) & x(61) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(79) & x(82) & x(83) & x(84) & x(85) & x(87) & x(88) & x(90) & x(91) & x(92) & x(93) & x(94) & x(95) & x(96) & x(101) & x(102) & x(103) & x(104) & x(105) & x(106) & x(107) & x(108) & x(110) & x(111) & x(112) & x(113) & x(115) & x(139) & x(140) & x(141) & x(142) & x(167) & x(168) & x(169) & x(196) & x(220) & x(221) & x(222) & x(248) & x(249) & x(250) & x(276) & x(277) & x(278) & x(305) & x(306) & x(333) & x(348) & x(349) & x(350) & x(364) & x(367) & x(378) & x(379) & x(392) & x(396) & x(397) & x(401) & x(406) & x(417) & x(419) & x(420) & x(422) & x(424) & x(425) & x(426) & x(427) & x(445) & x(448) & x(449) & x(450) & x(451) & x(453) & x(456) & x(476) & x(478) & x(479) & x(482) & x(483) & x(484) & x(491) & x(503) & x(504) & x(507) & x(511) & x(512) & x(532) & x(534) & x(535) & x(560) & x(562) & x(563) & x(587) & x(588) & x(591) & x(615) & x(616) & x(617) & x(619) & x(620) & x(643) & x(644) & x(645) & x(647) & x(648) & x(653) & x(654) & x(659) & x(671) & x(672) & x(673) & x(674) & x(676) & x(679) & x(684) & x(685) & x(698) & x(699) & x(700) & x(701) & x(702) & x(725) & x(726) & x(727) & x(728) & x(729) & x(730) & x(731) & x(752) & x(753) & x(754) & x(755) & x(756) & x(757) & x(758) & x(759) & x(760) & x(767) & x(768) & x(769) & x(771) & x(774) & x(779) & x(780) & x(781) & x(782) & x(783);
    y(244) <= not(p244_out);
    p244 : perceptron
        Generic map (
            WEIGHTS => "11111111111111111111111111111111000000000000011111111100000000000000000011111100000000000000011111111111110000000000000001000111100110111101100111001111110111001001101110011100000111000001111111111111111111110000011111",
            SHIFT => 4,
            B => 544,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p244_in,
            y(0) => p244_out,
            y(1 to 17 - 1) => dummy244
        );


    p245_in <= x(34) & x(35) & x(36) & x(37) & x(38) & x(39) & x(40) & x(41) & x(42) & x(43) & x(45) & x(46) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(79) & x(90) & x(91) & x(92) & x(104) & x(105) & x(109) & x(146) & x(165) & x(166) & x(172) & x(173) & x(174) & x(193) & x(198) & x(199) & x(200) & x(202) & x(220) & x(221) & x(222) & x(227) & x(228) & x(247) & x(248) & x(249) & x(250) & x(269) & x(275) & x(276) & x(277) & x(280) & x(295) & x(296) & x(297) & x(298) & x(299) & x(311) & x(320) & x(323) & x(324) & x(325) & x(326) & x(348) & x(349) & x(359) & x(388) & x(418) & x(425) & x(426) & x(444) & x(446) & x(453) & x(473) & x(474) & x(475) & x(487) & x(501) & x(502) & x(529) & x(530) & x(531) & x(535) & x(542) & x(543) & x(557) & x(558) & x(584) & x(585) & x(619) & x(695) & x(706) & x(707) & x(708) & x(719) & x(720) & x(721) & x(722) & x(723) & x(735) & x(736) & x(737) & x(744) & x(749) & x(764) & x(769) & x(770) & x(772) & x(773) & x(774);
    y(245) <= not(p245_out);
    p245 : perceptron
        Generic map (
            WEIGHTS => "00000000000000000000000000000000000110011101111000110000100011111110111100001110111110111111001111101110000011110111111",
            SHIFT => 4,
            B => -181,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p245_in,
            y(0) => p245_out,
            y(1 to 17 - 1) => dummy245
        );


    p246_in <= x(35) & x(36) & x(37) & x(38) & x(39) & x(40) & x(41) & x(42) & x(46) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(79) & x(90) & x(91) & x(95) & x(96) & x(97) & x(98) & x(99) & x(100) & x(101) & x(102) & x(103) & x(104) & x(105) & x(106) & x(136) & x(164) & x(165) & x(192) & x(193) & x(198) & x(226) & x(280) & x(302) & x(307) & x(314) & x(315) & x(334) & x(353) & x(359) & x(361) & x(362) & x(379) & x(381) & x(385) & x(386) & x(387) & x(388) & x(390) & x(394) & x(401) & x(409) & x(413) & x(414) & x(415) & x(416) & x(418) & x(430) & x(446) & x(458) & x(475) & x(485) & x(509) & x(511) & x(543) & x(544) & x(553) & x(573) & x(584) & x(592) & x(612) & x(648) & x(657) & x(691) & x(719) & x(720) & x(736) & x(737) & x(750) & x(770) & x(773) & x(774);
    y(246) <= not(p246_out);
    p246 : perceptron
        Generic map (
            WEIGHTS => "11111111111111111111111111111111111111111000000000000001000011110010111101010111111111110000000000",
            SHIFT => 4,
            B => 473,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p246_in,
            y(0) => p246_out,
            y(1 to 16 - 1) => dummy246
        );


    p247_in <= x(37) & x(66) & x(68) & x(118) & x(133) & x(182) & x(183) & x(192) & x(211) & x(302) & x(303) & x(304) & x(306) & x(329) & x(330) & x(331) & x(332) & x(333) & x(361) & x(362) & x(386) & x(387) & x(389) & x(390) & x(414) & x(415) & x(416) & x(418) & x(445) & x(446) & x(447) & x(450) & x(473) & x(474) & x(475) & x(479) & x(501) & x(502) & x(507) & x(529) & x(535) & x(557) & x(563) & x(584) & x(591) & x(612) & x(619) & x(647) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(723) & x(744) & x(745) & x(746) & x(747) & x(748) & x(749);
    y(247) <= not(p247_out);
    p247 : perceptron
        Generic map (
            WEIGHTS => "1110100100000000000011001110000000000000000000000000000000000",
            SHIFT => 5,
            B => -1626,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p247_in,
            y(0) => p247_out,
            y(1 to 17 - 1) => dummy247
        );


    p248_in <= x(37) & x(45) & x(62) & x(63) & x(64) & x(65) & x(66) & x(68) & x(69) & x(70) & x(71) & x(72) & x(74) & x(75) & x(108) & x(118) & x(123) & x(124) & x(133) & x(134) & x(135) & x(136) & x(146) & x(151) & x(162) & x(164) & x(165) & x(172) & x(173) & x(174) & x(175) & x(176) & x(177) & x(192) & x(193) & x(194) & x(197) & x(200) & x(220) & x(221) & x(222) & x(242) & x(248) & x(249) & x(250) & x(276) & x(277) & x(296) & x(297) & x(298) & x(299) & x(300) & x(301) & x(302) & x(305) & x(309) & x(315) & x(316) & x(330) & x(331) & x(332) & x(338) & x(342) & x(350) & x(360) & x(361) & x(362) & x(366) & x(368) & x(377) & x(378) & x(390) & x(405) & x(422) & x(425) & x(434) & x(446) & x(450) & x(453) & x(455) & x(466) & x(473) & x(474) & x(479) & x(481) & x(489) & x(501) & x(502) & x(507) & x(529) & x(534) & x(535) & x(543) & x(544) & x(557) & x(558) & x(563) & x(564) & x(577) & x(581) & x(584) & x(591) & x(592) & x(612) & x(619) & x(647) & x(675) & x(692) & x(693) & x(694) & x(695) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(747) & x(748);
    y(248) <= not(p248_out);
    p248 : perceptron
        Generic map (
            WEIGHTS => "00000000000000111100001100011111100011000100000111111101001111001111000101101111111110111111001111111111111000000000000",
            SHIFT => 4,
            B => 60,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p248_in,
            y(0) => p248_out,
            y(1 to 17 - 1) => dummy248
        );


    p249_in <= x(40) & x(41) & x(63) & x(67) & x(68) & x(69) & x(70) & x(72) & x(76) & x(78) & x(79) & x(101) & x(102) & x(103) & x(104) & x(105) & x(106) & x(108) & x(165) & x(166) & x(171) & x(172) & x(191) & x(192) & x(193) & x(197) & x(200) & x(219) & x(220) & x(221) & x(226) & x(247) & x(248) & x(249) & x(250) & x(254) & x(275) & x(276) & x(277) & x(289) & x(290) & x(291) & x(295) & x(317) & x(330) & x(331) & x(332) & x(334) & x(358) & x(359) & x(360) & x(386) & x(414) & x(441) & x(450) & x(461) & x(467) & x(469) & x(478) & x(495) & x(506) & x(507) & x(534) & x(535) & x(549) & x(550) & x(562) & x(563) & x(577) & x(591) & x(618) & x(619) & x(620) & x(646) & x(647) & x(648) & x(665) & x(675) & x(676) & x(677) & x(678) & x(679);
    y(249) <= not(p249_out);
    p249 : perceptron
        Generic map (
            WEIGHTS => "0000000000000000001100111001111111111111110100010000000100000000000000000000100000",
            SHIFT => 4,
            B => -753,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p249_in,
            y(0) => p249_out,
            y(1 to 16 - 1) => dummy249
        );


    p250_in <= x(35) & x(37) & x(38) & x(40) & x(44) & x(45) & x(46) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(92) & x(93) & x(94) & x(107) & x(108) & x(163) & x(192) & x(193) & x(194) & x(198) & x(219) & x(220) & x(221) & x(222) & x(228) & x(248) & x(249) & x(250) & x(276) & x(277) & x(278) & x(297) & x(298) & x(299) & x(302) & x(303) & x(305) & x(306) & x(309) & x(310) & x(311) & x(326) & x(327) & x(328) & x(329) & x(330) & x(331) & x(332) & x(333) & x(337) & x(338) & x(346) & x(347) & x(348) & x(349) & x(350) & x(357) & x(358) & x(359) & x(360) & x(366) & x(373) & x(374) & x(375) & x(376) & x(377) & x(378) & x(394) & x(425) & x(453) & x(454) & x(479) & x(484) & x(485) & x(486) & x(489) & x(494) & x(501) & x(507) & x(512) & x(513) & x(514) & x(515) & x(517) & x(535) & x(545) & x(550) & x(557) & x(563) & x(591) & x(648) & x(649) & x(654) & x(655) & x(656) & x(677) & x(694) & x(720) & x(721) & x(723) & x(735) & x(736) & x(742) & x(743) & x(769) & x(770) & x(772) & x(773) & x(774);
    y(250) <= not(p250_out);
    p250 : perceptron
        Generic map (
            WEIGHTS => "11111111111111111111111001111011110111111000001100000000001001111100000111111000010000101000001010111111111111000000000",
            SHIFT => 4,
            B => 232,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p250_in,
            y(0) => p250_out,
            y(1 to 17 - 1) => dummy250
        );


    p251_in <= x(38) & x(39) & x(40) & x(41) & x(44) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(78) & x(79) & x(90) & x(91) & x(92) & x(93) & x(94) & x(95) & x(96) & x(100) & x(101) & x(102) & x(103) & x(104) & x(105) & x(136) & x(145) & x(172) & x(192) & x(193) & x(220) & x(221) & x(247) & x(248) & x(249) & x(250) & x(276) & x(277) & x(307) & x(310) & x(319) & x(320) & x(321) & x(322) & x(333) & x(334) & x(338) & x(339) & x(347) & x(348) & x(349) & x(350) & x(351) & x(361) & x(362) & x(366) & x(375) & x(376) & x(377) & x(378) & x(450) & x(473) & x(501) & x(502) & x(507) & x(517) & x(528) & x(529) & x(535) & x(542) & x(543) & x(544) & x(545) & x(556) & x(557) & x(571) & x(572) & x(584) & x(591) & x(611) & x(612) & x(638) & x(655) & x(656) & x(657) & x(658) & x(675) & x(690) & x(692) & x(693) & x(694) & x(695) & x(697) & x(719) & x(720) & x(721) & x(722) & x(741) & x(742) & x(743) & x(748) & x(764);
    y(251) <= not(p251_out);
    p251 : perceptron
        Generic map (
            WEIGHTS => "11111111111111111111111111111100000000000000100000011000000010000011101110111111111011100000000001000011101",
            SHIFT => 4,
            B => 161,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p251_in,
            y(0) => p251_out,
            y(1 to 16 - 1) => dummy251
        );


    p252_in <= x(35) & x(63) & x(68) & x(108) & x(164) & x(165) & x(177) & x(178) & x(191) & x(192) & x(193) & x(197) & x(198) & x(220) & x(221) & x(226) & x(247) & x(248) & x(249) & x(250) & x(254) & x(266) & x(276) & x(277) & x(282) & x(292) & x(294) & x(305) & x(309) & x(310) & x(329) & x(330) & x(331) & x(338) & x(339) & x(347) & x(348) & x(357) & x(358) & x(366) & x(367) & x(374) & x(375) & x(376) & x(394) & x(397) & x(400) & x(416) & x(424) & x(425) & x(444) & x(445) & x(450) & x(472) & x(490) & x(494) & x(515) & x(516) & x(524) & x(534) & x(535) & x(544) & x(550) & x(578) & x(592) & x(618) & x(620) & x(621) & x(647) & x(674) & x(675) & x(677) & x(682) & x(703) & x(711) & x(714) & x(715) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(736) & x(737) & x(738) & x(739) & x(740) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(750) & x(764) & x(765) & x(766) & x(769) & x(770) & x(771) & x(772) & x(773) & x(774);
    y(252) <= not(p252_out);
    p252 : perceptron
        Generic map (
            WEIGHTS => "0000111111110110111100110001000000011000011101111110110100111011111111111100000000000000000000000000000000",
            SHIFT => 4,
            B => -275,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p252_in,
            y(0) => p252_out,
            y(1 to 16 - 1) => dummy252
        );


    p253_in <= x(37) & x(38) & x(39) & x(40) & x(41) & x(45) & x(46) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(79) & x(99) & x(100) & x(102) & x(103) & x(104) & x(105) & x(106) & x(133) & x(135) & x(163) & x(164) & x(165) & x(182) & x(183) & x(184) & x(191) & x(192) & x(193) & x(194) & x(210) & x(211) & x(212) & x(219) & x(220) & x(221) & x(222) & x(227) & x(238) & x(239) & x(247) & x(248) & x(249) & x(250) & x(254) & x(276) & x(277) & x(283) & x(301) & x(302) & x(303) & x(304) & x(310) & x(311) & x(312) & x(320) & x(327) & x(328) & x(329) & x(330) & x(331) & x(332) & x(339) & x(347) & x(348) & x(357) & x(358) & x(359) & x(360) & x(361) & x(390) & x(414) & x(418) & x(425) & x(446) & x(453) & x(454) & x(473) & x(474) & x(475) & x(481) & x(501) & x(502) & x(514) & x(529) & x(557) & x(558) & x(619) & x(675) & x(677) & x(678) & x(679) & x(695) & x(704) & x(705) & x(706) & x(707) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(732) & x(735) & x(747) & x(748) & x(749) & x(761) & x(769) & x(770) & x(771) & x(773);
    y(253) <= not(p253_out);
    p253 : perceptron
        Generic map (
            WEIGHTS => "111111111111111111111111111111111111100011110001111100111111110000111100000011100000010000000000000000111101111000000000100011111",
            SHIFT => 4,
            B => 560,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p253_in,
            y(0) => p253_out,
            y(1 to 17 - 1) => dummy253
        );


    p254_in <= x(37) & x(38) & x(39) & x(40) & x(41) & x(62) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(79) & x(99) & x(100) & x(103) & x(104) & x(105) & x(106) & x(198) & x(199) & x(201) & x(202) & x(204) & x(210) & x(211) & x(218) & x(226) & x(227) & x(228) & x(229) & x(254) & x(255) & x(256) & x(257) & x(268) & x(269) & x(270) & x(271) & x(280) & x(281) & x(282) & x(283) & x(284) & x(285) & x(296) & x(297) & x(307) & x(309) & x(310) & x(311) & x(312) & x(337) & x(338) & x(339) & x(350) & x(361) & x(362) & x(366) & x(367) & x(377) & x(378) & x(379) & x(381) & x(382) & x(386) & x(389) & x(390) & x(394) & x(405) & x(418) & x(446) & x(453) & x(454) & x(473) & x(474) & x(481) & x(482) & x(487) & x(500) & x(501) & x(502) & x(514) & x(515) & x(528) & x(529) & x(556) & x(557) & x(584) & x(692) & x(693) & x(694) & x(695) & x(696) & x(706) & x(707) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(735) & x(736) & x(743) & x(748) & x(749) & x(761) & x(764) & x(765) & x(766) & x(769) & x(770) & x(771) & x(772) & x(773) & x(774);
    y(254) <= not(p254_out);
    p254 : perceptron
        Generic map (
            WEIGHTS => "0000000000000000000000000000011111001111111111111111111111111111101111000000111011111111011100111110000011000000111001111111111",
            SHIFT => 4,
            B => 392,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p254_in,
            y(0) => p254_out,
            y(1 to 17 - 1) => dummy254
        );


    p255_in <= x(35) & x(63) & x(66) & x(67) & x(68) & x(69) & x(91) & x(108) & x(135) & x(163) & x(164) & x(182) & x(183) & x(191) & x(192) & x(197) & x(210) & x(211) & x(212) & x(220) & x(221) & x(237) & x(238) & x(239) & x(248) & x(249) & x(266) & x(277) & x(283) & x(301) & x(302) & x(303) & x(304) & x(328) & x(329) & x(330) & x(331) & x(332) & x(347) & x(350) & x(356) & x(357) & x(358) & x(359) & x(397) & x(400) & x(450) & x(487) & x(507) & x(513) & x(514) & x(515) & x(516) & x(535) & x(542) & x(543) & x(563) & x(591) & x(647) & x(648) & x(675) & x(676) & x(677) & x(678) & x(691) & x(692) & x(695) & x(703) & x(705) & x(706) & x(708) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(735) & x(739) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(748) & x(749);
    y(255) <= not(p255_out);
    p255 : perceptron
        Generic map (
            WEIGHTS => "111111110001100011100111001001111111110111110001011110110000000011100001111111101111111111",
            SHIFT => 4,
            B => 206,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p255_in,
            y(0) => p255_out,
            y(1 to 16 - 1) => dummy255
        );



--    p1 : perceptron
--        Generic map (
--            WEIGHTS => "",
--            SHIFT => "",
--            B => "",
--            BATCH_POSITIVE => ""
--        )
--        Port map (
--            x => x(0) & x(2) & ...,
--            y => ""
--        );

end layer_1;

architecture layer_2 of layer is

    Component perceptron
    Generic (
        WEIGHTS : STD_LOGIC_VECTOR := (others => '0');
        SHIFT : Integer;     -- number of shift (left + or right -)
        B : Integer;          -- bias of batch norm
        BATCH_POSITIVE : Boolean    
    );
    Port ( 
        x : in STD_LOGIC_VECTOR;
        y : out STD_LOGIC_VECTOR
   );
    end component;
    
    -- Signals
    signal p0_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p0_out : STD_LOGIC;
	signal p1_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p1_out : STD_LOGIC;
	signal p2_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p2_out : STD_LOGIC;
	signal p3_in : STD_LOGIC_VECTOR(0 to 10 - 1);
	signal p3_out : STD_LOGIC;
	signal p4_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p4_out : STD_LOGIC;
	signal p5_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p5_out : STD_LOGIC;
	signal p6_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p6_out : STD_LOGIC;
	signal p7_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p7_out : STD_LOGIC;
	signal p8_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p8_out : STD_LOGIC;
	signal p9_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p9_out : STD_LOGIC;
	signal p10_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p10_out : STD_LOGIC;
	signal p11_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p11_out : STD_LOGIC;
	signal p12_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p12_out : STD_LOGIC;
	signal p13_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p13_out : STD_LOGIC;
	signal p14_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p14_out : STD_LOGIC;
	signal p15_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p15_out : STD_LOGIC;
	signal p16_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p16_out : STD_LOGIC;
	signal p17_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p17_out : STD_LOGIC;
	signal p18_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p18_out : STD_LOGIC;
	signal p19_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p19_out : STD_LOGIC;
	signal p20_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p20_out : STD_LOGIC;
	signal p21_in : STD_LOGIC_VECTOR(0 to 7 - 1);
	signal p21_out : STD_LOGIC;
	signal p22_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p22_out : STD_LOGIC;
	signal p23_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p23_out : STD_LOGIC;
	signal p24_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p24_out : STD_LOGIC;
	signal p25_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p25_out : STD_LOGIC;
	signal p26_in : STD_LOGIC_VECTOR(0 to 8 - 1);
	signal p26_out : STD_LOGIC;
	signal p27_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p27_out : STD_LOGIC;
	signal p28_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p28_out : STD_LOGIC;
	signal p29_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p29_out : STD_LOGIC;
	signal p30_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p30_out : STD_LOGIC;
	signal p31_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p31_out : STD_LOGIC;
	signal p32_in : STD_LOGIC_VECTOR(0 to 7 - 1);
	signal p32_out : STD_LOGIC;
	signal p33_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p33_out : STD_LOGIC;
	signal p34_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p34_out : STD_LOGIC;
	signal p35_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p35_out : STD_LOGIC;
	signal p36_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p36_out : STD_LOGIC;
	signal p37_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p37_out : STD_LOGIC;
	signal p38_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p38_out : STD_LOGIC;
	signal p39_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p39_out : STD_LOGIC;
	signal p40_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p40_out : STD_LOGIC;
	signal p41_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p41_out : STD_LOGIC;
	signal p42_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p42_out : STD_LOGIC;
	signal p43_in : STD_LOGIC_VECTOR(0 to 7 - 1);
	signal p43_out : STD_LOGIC;
	signal p44_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p44_out : STD_LOGIC;
	signal p45_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p45_out : STD_LOGIC;
	signal p46_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p46_out : STD_LOGIC;
	signal p47_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p47_out : STD_LOGIC;
	signal p48_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p48_out : STD_LOGIC;
	signal p49_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p49_out : STD_LOGIC;
	signal p50_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p50_out : STD_LOGIC;
	signal p51_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p51_out : STD_LOGIC;
	signal p52_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p52_out : STD_LOGIC;
	signal p53_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p53_out : STD_LOGIC;
	signal p54_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p54_out : STD_LOGIC;
	signal p55_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p55_out : STD_LOGIC;
	signal p56_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p56_out : STD_LOGIC;
	signal p57_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p57_out : STD_LOGIC;
	signal p58_in : STD_LOGIC_VECTOR(0 to 7 - 1);
	signal p58_out : STD_LOGIC;
	signal p59_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p59_out : STD_LOGIC;
	signal p60_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p60_out : STD_LOGIC;
	signal p61_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p61_out : STD_LOGIC;
	signal p62_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p62_out : STD_LOGIC;
	signal p63_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p63_out : STD_LOGIC;
	signal p64_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p64_out : STD_LOGIC;
	signal p65_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p65_out : STD_LOGIC;
	signal p66_in : STD_LOGIC_VECTOR(0 to 7 - 1);
	signal p66_out : STD_LOGIC;
	signal p67_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p67_out : STD_LOGIC;
	signal p68_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p68_out : STD_LOGIC;
	signal p69_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p69_out : STD_LOGIC;
	signal p70_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p70_out : STD_LOGIC;
	signal p71_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p71_out : STD_LOGIC;
	signal p72_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p72_out : STD_LOGIC;
	signal p73_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p73_out : STD_LOGIC;
	signal p74_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p74_out : STD_LOGIC;
	signal p75_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p75_out : STD_LOGIC;
	signal p76_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p76_out : STD_LOGIC;
	signal p77_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p77_out : STD_LOGIC;
	signal p78_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p78_out : STD_LOGIC;
	signal p79_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p79_out : STD_LOGIC;
	signal p80_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p80_out : STD_LOGIC;
	signal p81_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p81_out : STD_LOGIC;
	signal p82_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p82_out : STD_LOGIC;
	signal p83_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p83_out : STD_LOGIC;
	signal p84_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p84_out : STD_LOGIC;
	signal p85_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p85_out : STD_LOGIC;
	signal p86_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p86_out : STD_LOGIC;
	signal p87_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p87_out : STD_LOGIC;
	signal p88_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p88_out : STD_LOGIC;
	signal p89_in : STD_LOGIC_VECTOR(0 to 7 - 1);
	signal p89_out : STD_LOGIC;
	signal p90_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p90_out : STD_LOGIC;
	signal p91_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p91_out : STD_LOGIC;
	signal p92_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p92_out : STD_LOGIC;
	signal p93_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p93_out : STD_LOGIC;
	signal p94_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p94_out : STD_LOGIC;
	signal p95_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p95_out : STD_LOGIC;
	signal p96_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p96_out : STD_LOGIC;
	signal p97_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p97_out : STD_LOGIC;
	signal p98_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p98_out : STD_LOGIC;
	signal p99_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p99_out : STD_LOGIC;
	signal p100_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p100_out : STD_LOGIC;
	signal p101_in : STD_LOGIC_VECTOR(0 to 7 - 1);
	signal p101_out : STD_LOGIC;
	signal p102_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p102_out : STD_LOGIC;
	signal p103_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p103_out : STD_LOGIC;
	signal p104_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p104_out : STD_LOGIC;
	signal p105_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p105_out : STD_LOGIC;
	signal p106_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p106_out : STD_LOGIC;
	signal p107_in : STD_LOGIC_VECTOR(0 to 10 - 1);
	signal p107_out : STD_LOGIC;
	signal p108_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p108_out : STD_LOGIC;
	signal p109_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p109_out : STD_LOGIC;
	signal p110_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p110_out : STD_LOGIC;
	signal p111_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p111_out : STD_LOGIC;
	signal p112_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p112_out : STD_LOGIC;
	signal p113_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p113_out : STD_LOGIC;
	signal p114_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p114_out : STD_LOGIC;
	signal p115_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p115_out : STD_LOGIC;
	signal p116_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p116_out : STD_LOGIC;
	signal p117_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p117_out : STD_LOGIC;
	signal p118_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p118_out : STD_LOGIC;
	signal p119_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p119_out : STD_LOGIC;
	signal p120_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p120_out : STD_LOGIC;
	signal p121_in : STD_LOGIC_VECTOR(0 to 9 - 1);
	signal p121_out : STD_LOGIC;
	signal p122_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p122_out : STD_LOGIC;
	signal p123_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p123_out : STD_LOGIC;
	signal p124_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p124_out : STD_LOGIC;
	signal p125_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p125_out : STD_LOGIC;
	signal p126_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p126_out : STD_LOGIC;
	signal p127_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p127_out : STD_LOGIC;
	signal p128_in : STD_LOGIC_VECTOR(0 to 7 - 1);
	signal p128_out : STD_LOGIC;
	signal p129_in : STD_LOGIC_VECTOR(0 to 8 - 1);
	signal p129_out : STD_LOGIC;
	signal p130_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p130_out : STD_LOGIC;
	signal p131_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p131_out : STD_LOGIC;
	signal p132_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p132_out : STD_LOGIC;
	signal p133_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p133_out : STD_LOGIC;
	signal p134_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p134_out : STD_LOGIC;
	signal p135_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p135_out : STD_LOGIC;
	signal p136_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p136_out : STD_LOGIC;
	signal p137_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p137_out : STD_LOGIC;
	signal p138_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p138_out : STD_LOGIC;
	signal p139_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p139_out : STD_LOGIC;
	signal p140_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p140_out : STD_LOGIC;
	signal p141_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p141_out : STD_LOGIC;
	signal p142_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p142_out : STD_LOGIC;
	signal p143_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p143_out : STD_LOGIC;
	signal p144_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p144_out : STD_LOGIC;
	signal p145_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p145_out : STD_LOGIC;
	signal p146_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p146_out : STD_LOGIC;
	signal p147_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p147_out : STD_LOGIC;
	signal p148_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p148_out : STD_LOGIC;
	signal p149_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p149_out : STD_LOGIC;
	signal p150_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p150_out : STD_LOGIC;
	signal p151_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p151_out : STD_LOGIC;
	signal p152_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p152_out : STD_LOGIC;
	signal p153_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p153_out : STD_LOGIC;
	signal p154_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p154_out : STD_LOGIC;
	signal p155_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p155_out : STD_LOGIC;
	signal p156_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p156_out : STD_LOGIC;
	signal p157_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p157_out : STD_LOGIC;
	signal p159_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p159_out : STD_LOGIC;
	signal p160_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p160_out : STD_LOGIC;
	signal p161_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p161_out : STD_LOGIC;
	signal p162_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p162_out : STD_LOGIC;
	signal p163_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p163_out : STD_LOGIC;
	signal p164_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p164_out : STD_LOGIC;
	signal p165_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p165_out : STD_LOGIC;
	signal p166_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p166_out : STD_LOGIC;
	signal p167_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p167_out : STD_LOGIC;
	signal p168_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p168_out : STD_LOGIC;
	signal p169_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p169_out : STD_LOGIC;
	signal p170_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p170_out : STD_LOGIC;
	signal p171_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p171_out : STD_LOGIC;
	signal p172_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p172_out : STD_LOGIC;
	signal p173_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p173_out : STD_LOGIC;
	signal p174_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p174_out : STD_LOGIC;
	signal p175_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p175_out : STD_LOGIC;
	signal p176_in : STD_LOGIC_VECTOR(0 to 7 - 1);
	signal p176_out : STD_LOGIC;
	signal p177_in : STD_LOGIC_VECTOR(0 to 7 - 1);
	signal p177_out : STD_LOGIC;
	signal p178_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p178_out : STD_LOGIC;
	signal p179_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p179_out : STD_LOGIC;
	signal p180_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p180_out : STD_LOGIC;
	signal p181_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p181_out : STD_LOGIC;
	signal p182_in : STD_LOGIC_VECTOR(0 to 9 - 1);
	signal p182_out : STD_LOGIC;
	signal p183_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p183_out : STD_LOGIC;
	signal p184_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p184_out : STD_LOGIC;
	signal p185_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p185_out : STD_LOGIC;
	signal p186_in : STD_LOGIC_VECTOR(0 to 8 - 1);
	signal p186_out : STD_LOGIC;
	signal p187_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p187_out : STD_LOGIC;
	signal p188_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p188_out : STD_LOGIC;
	signal p189_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p189_out : STD_LOGIC;
	signal p190_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p190_out : STD_LOGIC;
	signal p191_in : STD_LOGIC_VECTOR(0 to 7 - 1);
	signal p191_out : STD_LOGIC;
	signal p192_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p192_out : STD_LOGIC;
	signal p193_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p193_out : STD_LOGIC;
	signal p194_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p194_out : STD_LOGIC;
	signal p195_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p195_out : STD_LOGIC;
	signal p196_in : STD_LOGIC_VECTOR(0 to 7 - 1);
	signal p196_out : STD_LOGIC;
	signal p197_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p197_out : STD_LOGIC;
	signal p198_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p198_out : STD_LOGIC;
	signal p199_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p199_out : STD_LOGIC;
	signal p200_in : STD_LOGIC_VECTOR(0 to 9 - 1);
	signal p200_out : STD_LOGIC;
	signal p201_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p201_out : STD_LOGIC;
	signal p202_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p202_out : STD_LOGIC;
	signal p203_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p203_out : STD_LOGIC;
	signal p204_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p204_out : STD_LOGIC;
	signal p205_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p205_out : STD_LOGIC;
	signal p206_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p206_out : STD_LOGIC;
	signal p207_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p207_out : STD_LOGIC;
	signal p208_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p208_out : STD_LOGIC;
	signal p209_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p209_out : STD_LOGIC;
	signal p210_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p210_out : STD_LOGIC;
	signal p211_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p211_out : STD_LOGIC;
	signal p212_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p212_out : STD_LOGIC;
	signal p213_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p213_out : STD_LOGIC;
	signal p214_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p214_out : STD_LOGIC;
	signal p215_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p215_out : STD_LOGIC;
	signal p216_in : STD_LOGIC_VECTOR(0 to 7 - 1);
	signal p216_out : STD_LOGIC;
	signal p217_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p217_out : STD_LOGIC;
	signal p218_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p218_out : STD_LOGIC;
	signal p219_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p219_out : STD_LOGIC;
	signal p220_in : STD_LOGIC_VECTOR(0 to 8 - 1);
	signal p220_out : STD_LOGIC;
	signal p221_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p221_out : STD_LOGIC;
	signal p222_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p222_out : STD_LOGIC;
	signal p223_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p223_out : STD_LOGIC;
	signal p224_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p224_out : STD_LOGIC;
	signal p225_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p225_out : STD_LOGIC;
	signal p226_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p226_out : STD_LOGIC;
	signal p227_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p227_out : STD_LOGIC;
	signal p228_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p228_out : STD_LOGIC;
	signal p229_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p229_out : STD_LOGIC;
	signal p230_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p230_out : STD_LOGIC;
	signal p231_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p231_out : STD_LOGIC;
	signal p232_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p232_out : STD_LOGIC;
	signal p233_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p233_out : STD_LOGIC;
	signal p234_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p234_out : STD_LOGIC;
	signal p235_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p235_out : STD_LOGIC;
	signal p236_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p236_out : STD_LOGIC;
	signal p237_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p237_out : STD_LOGIC;
	signal p238_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p238_out : STD_LOGIC;
	signal p239_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p239_out : STD_LOGIC;
	signal p240_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p240_out : STD_LOGIC;
	signal p241_in : STD_LOGIC_VECTOR(0 to 8 - 1);
	signal p241_out : STD_LOGIC;
	signal p242_in : STD_LOGIC_VECTOR(0 to 8 - 1);
	signal p242_out : STD_LOGIC;
	signal p243_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p243_out : STD_LOGIC;
	signal p244_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p244_out : STD_LOGIC;
	signal p245_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p245_out : STD_LOGIC;
	signal p246_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p246_out : STD_LOGIC;
	signal p247_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p247_out : STD_LOGIC;
	signal p248_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p248_out : STD_LOGIC;
	signal p249_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p249_out : STD_LOGIC;
	signal p250_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p250_out : STD_LOGIC;
	signal p251_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p251_out : STD_LOGIC;
	signal p252_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p252_out : STD_LOGIC;
	signal p253_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p253_out : STD_LOGIC;
	signal p254_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p254_out : STD_LOGIC;
	signal p255_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p255_out : STD_LOGIC;
	
    
    -- Dummies
    signal dummy0 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy1 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy2 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy3 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy4 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy5 : STD_LOGIC_VECTOR(0 to 11 - 2);
	signal dummy6 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy7 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy8 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy9 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy10 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy11 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy12 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy13 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy14 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy15 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy16 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy17 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy18 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy19 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy20 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy21 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy22 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy23 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy24 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy25 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy26 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy27 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy28 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy29 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy30 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy31 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy32 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy33 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy34 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy35 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy36 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy37 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy38 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy39 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy40 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy41 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy42 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy43 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy44 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy45 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy46 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy47 : STD_LOGIC_VECTOR(0 to 11 - 2);
	signal dummy48 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy49 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy50 : STD_LOGIC_VECTOR(0 to 11 - 2);
	signal dummy51 : STD_LOGIC_VECTOR(0 to 11 - 2);
	signal dummy52 : STD_LOGIC_VECTOR(0 to 11 - 2);
	signal dummy53 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy54 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy55 : STD_LOGIC_VECTOR(0 to 11 - 2);
	signal dummy56 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy57 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy58 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy59 : STD_LOGIC_VECTOR(0 to 11 - 2);
	signal dummy60 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy61 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy62 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy63 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy64 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy65 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy66 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy67 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy68 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy69 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy70 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy71 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy72 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy73 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy74 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy75 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy76 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy77 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy78 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy79 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy80 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy81 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy82 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy83 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy84 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy85 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy86 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy87 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy88 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy89 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy90 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy91 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy92 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy93 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy94 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy95 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy96 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy97 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy98 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy99 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy100 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy101 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy102 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy103 : STD_LOGIC_VECTOR(0 to 11 - 2);
	signal dummy104 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy105 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy106 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy107 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy108 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy109 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy110 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy111 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy112 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy113 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy114 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy115 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy116 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy117 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy118 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy119 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy120 : STD_LOGIC_VECTOR(0 to 11 - 2);
	signal dummy121 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy122 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy123 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy124 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy125 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy126 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy127 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy128 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy129 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy130 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy131 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy132 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy133 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy134 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy135 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy136 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy137 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy138 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy139 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy140 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy141 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy142 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy143 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy144 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy145 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy146 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy147 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy148 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy149 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy150 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy151 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy152 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy153 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy154 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy155 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy156 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy157 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy159 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy160 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy161 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy162 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy163 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy164 : STD_LOGIC_VECTOR(0 to 11 - 2);
	signal dummy165 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy166 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy167 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy168 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy169 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy170 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy171 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy172 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy173 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy174 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy175 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy176 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy177 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy178 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy179 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy180 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy181 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy182 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy183 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy184 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy185 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy186 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy187 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy188 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy189 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy190 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy191 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy192 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy193 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy194 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy195 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy196 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy197 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy198 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy199 : STD_LOGIC_VECTOR(0 to 11 - 2);
	signal dummy200 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy201 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy202 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy203 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy204 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy205 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy206 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy207 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy208 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy209 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy210 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy211 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy212 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy213 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy214 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy215 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy216 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy217 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy218 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy219 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy220 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy221 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy222 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy223 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy224 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy225 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy226 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy227 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy228 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy229 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy230 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy231 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy232 : STD_LOGIC_VECTOR(0 to 11 - 2);
	signal dummy233 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy234 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy235 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy236 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy237 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy238 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy239 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy240 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy241 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy242 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy243 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy244 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy245 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy246 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy247 : STD_LOGIC_VECTOR(0 to 11 - 2);
	signal dummy248 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy249 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy250 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy251 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy252 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy253 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy254 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy255 : STD_LOGIC_VECTOR(0 to 11 - 2);
	 
    
begin

    
    p0_in <= x(46) & x(79) & x(164) & x(188) & x(244);
    y(0) <= not(p0_out);
    p0 : perceptron
        Generic map (
            WEIGHTS => "10011",
            SHIFT => 5,
            B => 4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p0_in,
            y(0) => p0_out,
            y(1 to 13 - 1) => dummy0
        );


    p1_in <= x(18) & x(159);
    y(1) <= not(p1_out);
    p1 : perceptron
        Generic map (
            WEIGHTS => "01",
            SHIFT => 6,
            B => -8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p1_in,
            y(0) => p1_out,
            y(1 to 12 - 1) => dummy1
        );


    p2_in <= x(126) & x(152) & x(193) & x(244);
    y(2) <= not(p2_out);
    p2 : perceptron
        Generic map (
            WEIGHTS => "1000",
            SHIFT => 6,
            B => -12,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p2_in,
            y(0) => p2_out,
            y(1 to 14 - 1) => dummy2
        );


    p3_in <= x(48) & x(81) & x(93) & x(97) & x(99) & x(114) & x(122) & x(149) & x(188) & x(254);
    y(3) <= not(p3_out);
    p3 : perceptron
        Generic map (
            WEIGHTS => "0110010001",
            SHIFT => 4,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p3_in,
            y(0) => p3_out,
            y(1 to 13 - 1) => dummy3
        );


    p4_in <= x(56) & x(81) & x(128);
    y(4) <= not(p4_out);
    p4 : perceptron
        Generic map (
            WEIGHTS => "100",
            SHIFT => 6,
            B => 8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p4_in,
            y(0) => p4_out,
            y(1 to 13 - 1) => dummy4
        );


    p5_in <= x(18) & x(172);
    y(5) <= not(p5_out);
    p5 : perceptron
        Generic map (
            WEIGHTS => "00",
            SHIFT => 5,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p5_in,
            y(0) => p5_out,
            y(1 to 11 - 1) => dummy5
        );


    p6_in(0) <= x(200);
    y(6) <= not(p6_out);
    p6 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p6_in,
            y(0) => p6_out,
            y(1 to 12 - 1) => dummy6
        );


    p7_in <= x(31) & x(101) & x(122) & x(156) & x(164);
    y(7) <= not(p7_out);
    p7 : perceptron
        Generic map (
            WEIGHTS => "01101",
            SHIFT => 5,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p7_in,
            y(0) => p7_out,
            y(1 to 13 - 1) => dummy7
        );


    p8_in(0) <= x(63);
    y(8) <= not(p8_out);
    p8 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => 9,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p8_in,
            y(0) => p8_out,
            y(1 to 12 - 1) => dummy8
        );


    p9_in <= x(81) & x(122) & x(169);
    y(9) <= not(p9_out);
    p9 : perceptron
        Generic map (
            WEIGHTS => "100",
            SHIFT => 5,
            B => 13,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p9_in,
            y(0) => p9_out,
            y(1 to 12 - 1) => dummy9
        );


    p10_in <= x(26) & x(46) & x(200) & x(229);
    y(10) <= not(p10_out);
    p10 : perceptron
        Generic map (
            WEIGHTS => "1100",
            SHIFT => 5,
            B => -7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p10_in,
            y(0) => p10_out,
            y(1 to 12 - 1) => dummy10
        );


    p11_in <= x(82) & x(144) & x(244);
    y(11) <= not(p11_out);
    p11 : perceptron
        Generic map (
            WEIGHTS => "001",
            SHIFT => 5,
            B => 4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p11_in,
            y(0) => p11_out,
            y(1 to 12 - 1) => dummy11
        );


    p12_in <= x(56) & x(99) & x(117) & x(193) & x(254);
    y(12) <= not(p12_out);
    p12 : perceptron
        Generic map (
            WEIGHTS => "11011",
            SHIFT => 5,
            B => 15,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p12_in,
            y(0) => p12_out,
            y(1 to 13 - 1) => dummy12
        );


    p13_in <= x(14) & x(150) & x(193);
    y(13) <= not(p13_out);
    p13 : perceptron
        Generic map (
            WEIGHTS => "001",
            SHIFT => 6,
            B => -12,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p13_in,
            y(0) => p13_out,
            y(1 to 13 - 1) => dummy13
        );


    p14_in <= x(94) & x(99) & x(150);
    y(14) <= not(p14_out);
    p14 : perceptron
        Generic map (
            WEIGHTS => "010",
            SHIFT => 6,
            B => 4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p14_in,
            y(0) => p14_out,
            y(1 to 13 - 1) => dummy14
        );


    p15_in <= x(19) & x(25) & x(164);
    y(15) <= not(p15_out);
    p15 : perceptron
        Generic map (
            WEIGHTS => "110",
            SHIFT => 5,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p15_in,
            y(0) => p15_out,
            y(1 to 12 - 1) => dummy15
        );


    p16_in <= x(11) & x(48) & x(91) & x(202);
    y(16) <= not(p16_out);
    p16 : perceptron
        Generic map (
            WEIGHTS => "0011",
            SHIFT => 5,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p16_in,
            y(0) => p16_out,
            y(1 to 12 - 1) => dummy16
        );


    p17_in <= x(60) & x(133) & x(245);
    y(17) <= not(p17_out);
    p17 : perceptron
        Generic map (
            WEIGHTS => "010",
            SHIFT => 6,
            B => 6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p17_in,
            y(0) => p17_out,
            y(1 to 13 - 1) => dummy17
        );


    p18_in <= x(23) & x(135) & x(146);
    y(18) <= not(p18_out);
    p18 : perceptron
        Generic map (
            WEIGHTS => "000",
            SHIFT => 5,
            B => -16,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p18_in,
            y(0) => p18_out,
            y(1 to 12 - 1) => dummy18
        );


    p19_in <= x(133) & x(155);
    y(19) <= not(p19_out);
    p19 : perceptron
        Generic map (
            WEIGHTS => "10",
            SHIFT => 6,
            B => 15,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p19_in,
            y(0) => p19_out,
            y(1 to 12 - 1) => dummy19
        );


    p20_in(0) <= x(229);
    y(20) <= not(p20_out);
    p20 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => -9,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p20_in,
            y(0) => p20_out,
            y(1 to 12 - 1) => dummy20
        );


    p21_in <= x(104) & x(177) & x(188) & x(213) & x(224) & x(229) & x(239);
    y(21) <= not(p21_out);
    p21 : perceptron
        Generic map (
            WEIGHTS => "1000101",
            SHIFT => 5,
            B => -18,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p21_in,
            y(0) => p21_out,
            y(1 to 13 - 1) => dummy21
        );


    p22_in <= x(11) & x(26) & x(111) & x(116);
    y(22) <= not(p22_out);
    p22 : perceptron
        Generic map (
            WEIGHTS => "0110",
            SHIFT => 6,
            B => -15,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p22_in,
            y(0) => p22_out,
            y(1 to 13 - 1) => dummy22
        );


    p23_in(0) <= x(172);
    y(23) <= not(p23_out);
    p23 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p23_in,
            y(0) => p23_out,
            y(1 to 12 - 1) => dummy23
        );


    p24_in <= x(68) & x(81) & x(122) & x(133) & x(221);
    y(24) <= not(p24_out);
    p24 : perceptron
        Generic map (
            WEIGHTS => "11011",
            SHIFT => 5,
            B => 14,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p24_in,
            y(0) => p24_out,
            y(1 to 13 - 1) => dummy24
        );


    p25_in <= x(40) & x(51) & x(152);
    y(25) <= not(p25_out);
    p25 : perceptron
        Generic map (
            WEIGHTS => "100",
            SHIFT => 5,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p25_in,
            y(0) => p25_out,
            y(1 to 12 - 1) => dummy25
        );


    p26_in <= x(56) & x(99) & x(123) & x(152) & x(175) & x(193) & x(231) & x(254);
    y(26) <= not(p26_out);
    p26 : perceptron
        Generic map (
            WEIGHTS => "00011010",
            SHIFT => 4,
            B => -6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p26_in,
            y(0) => p26_out,
            y(1 to 13 - 1) => dummy26
        );


    p27_in <= x(152) & x(193) & x(200) & x(244);
    y(27) <= not(p27_out);
    p27 : perceptron
        Generic map (
            WEIGHTS => "0000",
            SHIFT => 6,
            B => -14,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p27_in,
            y(0) => p27_out,
            y(1 to 14 - 1) => dummy27
        );


    p28_in <= x(39) & x(193);
    y(28) <= not(p28_out);
    p28 : perceptron
        Generic map (
            WEIGHTS => "10",
            SHIFT => 6,
            B => -9,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p28_in,
            y(0) => p28_out,
            y(1 to 12 - 1) => dummy28
        );


    p29_in <= x(5) & x(60) & x(63) & x(105);
    y(29) <= not(p29_out);
    p29 : perceptron
        Generic map (
            WEIGHTS => "1000",
            SHIFT => 5,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p29_in,
            y(0) => p29_out,
            y(1 to 12 - 1) => dummy29
        );


    p30_in <= x(60) & x(134) & x(157) & x(193) & x(241);
    y(30) <= not(p30_out);
    p30 : perceptron
        Generic map (
            WEIGHTS => "00001",
            SHIFT => 5,
            B => -7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p30_in,
            y(0) => p30_out,
            y(1 to 13 - 1) => dummy30
        );


    p31_in <= x(48) & x(173);
    y(31) <= not(p31_out);
    p31 : perceptron
        Generic map (
            WEIGHTS => "10",
            SHIFT => 6,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p31_in,
            y(0) => p31_out,
            y(1 to 12 - 1) => dummy31
        );


    p32_in <= x(94) & x(117) & x(126) & x(150) & x(172) & x(193) & x(254);
    y(32) <= not(p32_out);
    p32 : perceptron
        Generic map (
            WEIGHTS => "1111100",
            SHIFT => 5,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p32_in,
            y(0) => p32_out,
            y(1 to 13 - 1) => dummy32
        );


    p33_in <= x(49) & x(222) & x(241);
    y(33) <= not(p33_out);
    p33 : perceptron
        Generic map (
            WEIGHTS => "010",
            SHIFT => 6,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p33_in,
            y(0) => p33_out,
            y(1 to 13 - 1) => dummy33
        );


    p34_in <= x(49) & x(54) & x(243);
    y(34) <= not(p34_out);
    p34 : perceptron
        Generic map (
            WEIGHTS => "011",
            SHIFT => 5,
            B => 8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p34_in,
            y(0) => p34_out,
            y(1 to 12 - 1) => dummy34
        );


    p35_in(0) <= x(202);
    y(35) <= not(p35_out);
    p35 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => -6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p35_in,
            y(0) => p35_out,
            y(1 to 12 - 1) => dummy35
        );


    p36_in <= x(40) & x(205) & x(225);
    y(36) <= not(p36_out);
    p36 : perceptron
        Generic map (
            WEIGHTS => "111",
            SHIFT => 5,
            B => 12,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p36_in,
            y(0) => p36_out,
            y(1 to 12 - 1) => dummy36
        );


    p37_in <= x(117) & x(142) & x(150) & x(157) & x(177);
    y(37) <= not(p37_out);
    p37 : perceptron
        Generic map (
            WEIGHTS => "11111",
            SHIFT => 5,
            B => 6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p37_in,
            y(0) => p37_out,
            y(1 to 13 - 1) => dummy37
        );


    p38_in <= x(69) & x(109) & x(231);
    y(38) <= not(p38_out);
    p38 : perceptron
        Generic map (
            WEIGHTS => "100",
            SHIFT => 5,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p38_in,
            y(0) => p38_out,
            y(1 to 12 - 1) => dummy38
        );


    p39_in <= x(40) & x(150);
    y(39) <= not(p39_out);
    p39 : perceptron
        Generic map (
            WEIGHTS => "10",
            SHIFT => 6,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p39_in,
            y(0) => p39_out,
            y(1 to 12 - 1) => dummy39
        );


    p40_in <= x(19) & x(142) & x(188);
    y(40) <= not(p40_out);
    p40 : perceptron
        Generic map (
            WEIGHTS => "000",
            SHIFT => 6,
            B => -24,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p40_in,
            y(0) => p40_out,
            y(1 to 13 - 1) => dummy40
        );


    p41_in <= x(39) & x(254);
    y(41) <= not(p41_out);
    p41 : perceptron
        Generic map (
            WEIGHTS => "01",
            SHIFT => 6,
            B => 16,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p41_in,
            y(0) => p41_out,
            y(1 to 12 - 1) => dummy41
        );


    p42_in <= x(200) & x(235) & x(254);
    y(42) <= not(p42_out);
    p42 : perceptron
        Generic map (
            WEIGHTS => "010",
            SHIFT => 6,
            B => -15,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p42_in,
            y(0) => p42_out,
            y(1 to 13 - 1) => dummy42
        );


    p43_in <= x(2) & x(126) & x(157) & x(177) & x(182) & x(239) & x(244);
    y(43) <= not(p43_out);
    p43 : perceptron
        Generic map (
            WEIGHTS => "1100011",
            SHIFT => 5,
            B => -20,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p43_in,
            y(0) => p43_out,
            y(1 to 13 - 1) => dummy43
        );


    p44_in <= x(132) & x(142) & x(188);
    y(44) <= not(p44_out);
    p44 : perceptron
        Generic map (
            WEIGHTS => "100",
            SHIFT => 5,
            B => -18,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p44_in,
            y(0) => p44_out,
            y(1 to 12 - 1) => dummy44
        );


    p45_in <= x(142) & x(172) & x(177) & x(188) & x(200) & x(229);
    y(45) <= not(p45_out);
    p45 : perceptron
        Generic map (
            WEIGHTS => "010000",
            SHIFT => 5,
            B => -15,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p45_in,
            y(0) => p45_out,
            y(1 to 13 - 1) => dummy45
        );


    p46_in <= x(101) & x(104);
    y(46) <= not(p46_out);
    p46 : perceptron
        Generic map (
            WEIGHTS => "10",
            SHIFT => 6,
            B => 13,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p46_in,
            y(0) => p46_out,
            y(1 to 12 - 1) => dummy46
        );


    p47_in(0) <= x(230);
    y(47) <= not(p47_out);
    p47 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 6,
            B => 10,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p47_in,
            y(0) => p47_out,
            y(1 to 11 - 1) => dummy47
        );


    p48_in <= x(119) & x(194);
    y(48) <= not(p48_out);
    p48 : perceptron
        Generic map (
            WEIGHTS => "00",
            SHIFT => 6,
            B => 7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p48_in,
            y(0) => p48_out,
            y(1 to 12 - 1) => dummy48
        );


    p49_in <= x(48) & x(68) & x(101) & x(122) & x(168) & x(169);
    y(49) <= not(p49_out);
    p49 : perceptron
        Generic map (
            WEIGHTS => "010000",
            SHIFT => 4,
            B => 18,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p49_in,
            y(0) => p49_out,
            y(1 to 12 - 1) => dummy49
        );


    p50_in <= x(15) & x(169);
    y(50) <= not(p50_out);
    p50 : perceptron
        Generic map (
            WEIGHTS => "11",
            SHIFT => 5,
            B => -15,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p50_in,
            y(0) => p50_out,
            y(1 to 11 - 1) => dummy50
        );


    p51_in(0) <= x(188);
    y(51) <= not(p51_out);
    p51 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 6,
            B => 8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p51_in,
            y(0) => p51_out,
            y(1 to 11 - 1) => dummy51
        );


    p52_in(0) <= x(183);
    y(52) <= not(p52_out);
    p52 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 6,
            B => -6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p52_in,
            y(0) => p52_out,
            y(1 to 11 - 1) => dummy52
        );


    p53_in <= x(60) & x(63) & x(165) & x(244);
    y(53) <= not(p53_out);
    p53 : perceptron
        Generic map (
            WEIGHTS => "0110",
            SHIFT => 5,
            B => -6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p53_in,
            y(0) => p53_out,
            y(1 to 12 - 1) => dummy53
        );


    p54_in <= x(99) & x(128) & x(231);
    y(54) <= not(p54_out);
    p54 : perceptron
        Generic map (
            WEIGHTS => "011",
            SHIFT => 5,
            B => -16,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p54_in,
            y(0) => p54_out,
            y(1 to 12 - 1) => dummy54
        );


    p55_in <= x(96) & x(104);
    y(55) <= not(p55_out);
    p55 : perceptron
        Generic map (
            WEIGHTS => "01",
            SHIFT => 5,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p55_in,
            y(0) => p55_out,
            y(1 to 11 - 1) => dummy55
        );


    p56_in <= x(195) & x(215) & x(248);
    y(56) <= not(p56_out);
    p56 : perceptron
        Generic map (
            WEIGHTS => "100",
            SHIFT => 6,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p56_in,
            y(0) => p56_out,
            y(1 to 13 - 1) => dummy56
        );


    p57_in <= x(35) & x(56) & x(144) & x(190) & x(203);
    y(57) <= not(p57_out);
    p57 : perceptron
        Generic map (
            WEIGHTS => "11001",
            SHIFT => 5,
            B => 6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p57_in,
            y(0) => p57_out,
            y(1 to 13 - 1) => dummy57
        );


    p58_in <= x(23) & x(99) & x(137) & x(152) & x(193) & x(200) & x(241);
    y(58) <= not(p58_out);
    p58 : perceptron
        Generic map (
            WEIGHTS => "1001110",
            SHIFT => 5,
            B => -10,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p58_in,
            y(0) => p58_out,
            y(1 to 13 - 1) => dummy58
        );


    p59_in <= x(116) & x(185);
    y(59) <= not(p59_out);
    p59 : perceptron
        Generic map (
            WEIGHTS => "00",
            SHIFT => 5,
            B => 9,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p59_in,
            y(0) => p59_out,
            y(1 to 11 - 1) => dummy59
        );


    p60_in <= x(63) & x(101) & x(122) & x(202);
    y(60) <= not(p60_out);
    p60 : perceptron
        Generic map (
            WEIGHTS => "1001",
            SHIFT => 5,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p60_in,
            y(0) => p60_out,
            y(1 to 13 - 1) => dummy60
        );


    p61_in(0) <= x(141);
    y(61) <= not(p61_out);
    p61 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p61_in,
            y(0) => p61_out,
            y(1 to 12 - 1) => dummy61
        );


    p62_in <= x(99) & x(175);
    y(62) <= not(p62_out);
    p62 : perceptron
        Generic map (
            WEIGHTS => "10",
            SHIFT => 6,
            B => 13,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p62_in,
            y(0) => p62_out,
            y(1 to 12 - 1) => dummy62
        );


    p63_in <= x(19) & x(208);
    y(63) <= not(p63_out);
    p63 : perceptron
        Generic map (
            WEIGHTS => "00",
            SHIFT => 6,
            B => -27,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p63_in,
            y(0) => p63_out,
            y(1 to 12 - 1) => dummy63
        );


    p64_in <= x(101) & x(172);
    y(64) <= not(p64_out);
    p64 : perceptron
        Generic map (
            WEIGHTS => "00",
            SHIFT => 6,
            B => -7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p64_in,
            y(0) => p64_out,
            y(1 to 12 - 1) => dummy64
        );


    p65_in <= x(51) & x(54) & x(133) & x(205);
    y(65) <= not(p65_out);
    p65 : perceptron
        Generic map (
            WEIGHTS => "1101",
            SHIFT => 6,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p65_in,
            y(0) => p65_out,
            y(1 to 13 - 1) => dummy65
        );


    p66_in <= x(8) & x(23) & x(109) & x(151) & x(200) & x(229) & x(235);
    y(66) <= not(p66_out);
    p66 : perceptron
        Generic map (
            WEIGHTS => "0110110",
            SHIFT => 5,
            B => 24,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p66_in,
            y(0) => p66_out,
            y(1 to 13 - 1) => dummy66
        );


    p67_in <= x(60) & x(63) & x(132) & x(144) & x(244);
    y(67) <= not(p67_out);
    p67 : perceptron
        Generic map (
            WEIGHTS => "01010",
            SHIFT => 5,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p67_in,
            y(0) => p67_out,
            y(1 to 13 - 1) => dummy67
        );


    p68_in <= x(12) & x(23) & x(200);
    y(68) <= not(p68_out);
    p68 : perceptron
        Generic map (
            WEIGHTS => "000",
            SHIFT => 5,
            B => -26,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p68_in,
            y(0) => p68_out,
            y(1 to 12 - 1) => dummy68
        );


    p69_in(0) <= x(37);
    y(69) <= not(p69_out);
    p69 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p69_in,
            y(0) => p69_out,
            y(1 to 12 - 1) => dummy69
        );


    p70_in <= x(37) & x(83) & x(164) & x(243);
    y(70) <= not(p70_out);
    p70 : perceptron
        Generic map (
            WEIGHTS => "1001",
            SHIFT => 5,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p70_in,
            y(0) => p70_out,
            y(1 to 12 - 1) => dummy70
        );


    p71_in <= x(48) & x(63);
    y(71) <= not(p71_out);
    p71 : perceptron
        Generic map (
            WEIGHTS => "00",
            SHIFT => 6,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p71_in,
            y(0) => p71_out,
            y(1 to 12 - 1) => dummy71
        );


    p72_in <= x(126) & x(150) & x(172) & x(193) & x(200) & x(229);
    y(72) <= not(p72_out);
    p72 : perceptron
        Generic map (
            WEIGHTS => "000111",
            SHIFT => 5,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p72_in,
            y(0) => p72_out,
            y(1 to 13 - 1) => dummy72
        );


    p73_in <= x(60) & x(152) & x(245);
    y(73) <= not(p73_out);
    p73 : perceptron
        Generic map (
            WEIGHTS => "000",
            SHIFT => 6,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p73_in,
            y(0) => p73_out,
            y(1 to 13 - 1) => dummy73
        );


    p74_in <= x(44) & x(63) & x(231) & x(243);
    y(74) <= not(p74_out);
    p74 : perceptron
        Generic map (
            WEIGHTS => "0100",
            SHIFT => 5,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p74_in,
            y(0) => p74_out,
            y(1 to 12 - 1) => dummy74
        );


    p75_in <= x(119) & x(202) & x(248);
    y(75) <= not(p75_out);
    p75 : perceptron
        Generic map (
            WEIGHTS => "100",
            SHIFT => 6,
            B => -12,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p75_in,
            y(0) => p75_out,
            y(1 to 13 - 1) => dummy75
        );


    p76_in <= x(91) & x(160) & x(243);
    y(76) <= not(p76_out);
    p76 : perceptron
        Generic map (
            WEIGHTS => "110",
            SHIFT => 5,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p76_in,
            y(0) => p76_out,
            y(1 to 12 - 1) => dummy76
        );


    p77_in <= x(97) & x(149);
    y(77) <= not(p77_out);
    p77 : perceptron
        Generic map (
            WEIGHTS => "00",
            SHIFT => 6,
            B => -11,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p77_in,
            y(0) => p77_out,
            y(1 to 12 - 1) => dummy77
        );


    p78_in <= x(39) & x(41) & x(79) & x(150);
    y(78) <= not(p78_out);
    p78 : perceptron
        Generic map (
            WEIGHTS => "0000",
            SHIFT => 5,
            B => 6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p78_in,
            y(0) => p78_out,
            y(1 to 12 - 1) => dummy78
        );


    p79_in <= x(9) & x(243);
    y(79) <= not(p79_out);
    p79 : perceptron
        Generic map (
            WEIGHTS => "00",
            SHIFT => 6,
            B => -10,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p79_in,
            y(0) => p79_out,
            y(1 to 12 - 1) => dummy79
        );


    p80_in <= x(39) & x(57) & x(58) & x(96) & x(99);
    y(80) <= not(p80_out);
    p80 : perceptron
        Generic map (
            WEIGHTS => "01000",
            SHIFT => 5,
            B => -14,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p80_in,
            y(0) => p80_out,
            y(1 to 13 - 1) => dummy80
        );


    p81_in <= x(63) & x(68) & x(231);
    y(81) <= not(p81_out);
    p81 : perceptron
        Generic map (
            WEIGHTS => "110",
            SHIFT => 6,
            B => -6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p81_in,
            y(0) => p81_out,
            y(1 to 13 - 1) => dummy81
        );


    p82_in(0) <= x(144);
    y(82) <= not(p82_out);
    p82 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p82_in,
            y(0) => p82_out,
            y(1 to 12 - 1) => dummy82
        );


    p83_in <= x(142) & x(150) & x(177);
    y(83) <= not(p83_out);
    p83 : perceptron
        Generic map (
            WEIGHTS => "000",
            SHIFT => 5,
            B => -15,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p83_in,
            y(0) => p83_out,
            y(1 to 12 - 1) => dummy83
        );


    p84_in <= x(128) & x(200) & x(240);
    y(84) <= not(p84_out);
    p84 : perceptron
        Generic map (
            WEIGHTS => "001",
            SHIFT => 6,
            B => 8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p84_in,
            y(0) => p84_out,
            y(1 to 13 - 1) => dummy84
        );


    p85_in <= x(56) & x(188);
    y(85) <= not(p85_out);
    p85 : perceptron
        Generic map (
            WEIGHTS => "11",
            SHIFT => 6,
            B => 8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p85_in,
            y(0) => p85_out,
            y(1 to 12 - 1) => dummy85
        );


    p86_in <= x(134) & x(144) & x(152) & x(164) & x(244);
    y(86) <= not(p86_out);
    p86 : perceptron
        Generic map (
            WEIGHTS => "01010",
            SHIFT => 5,
            B => -9,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p86_in,
            y(0) => p86_out,
            y(1 to 13 - 1) => dummy86
        );


    p87_in <= x(15) & x(38);
    y(87) <= not(p87_out);
    p87 : perceptron
        Generic map (
            WEIGHTS => "10",
            SHIFT => 6,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p87_in,
            y(0) => p87_out,
            y(1 to 12 - 1) => dummy87
        );


    p88_in(0) <= x(244);
    y(88) <= not(p88_out);
    p88 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => -18,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p88_in,
            y(0) => p88_out,
            y(1 to 12 - 1) => dummy88
        );


    p89_in <= x(63) & x(99) & x(111) & x(144) & x(152) & x(190) & x(254);
    y(89) <= not(p89_out);
    p89 : perceptron
        Generic map (
            WEIGHTS => "0000100",
            SHIFT => 5,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p89_in,
            y(0) => p89_out,
            y(1 to 13 - 1) => dummy89
        );


    p90_in <= x(81) & x(150) & x(152) & x(164) & x(252);
    y(90) <= not(p90_out);
    p90 : perceptron
        Generic map (
            WEIGHTS => "00010",
            SHIFT => 5,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p90_in,
            y(0) => p90_out,
            y(1 to 13 - 1) => dummy90
        );


    p91_in <= x(122) & x(231);
    y(91) <= not(p91_out);
    p91 : perceptron
        Generic map (
            WEIGHTS => "11",
            SHIFT => 6,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p91_in,
            y(0) => p91_out,
            y(1 to 12 - 1) => dummy91
        );


    p92_in <= x(5) & x(50);
    y(92) <= not(p92_out);
    p92 : perceptron
        Generic map (
            WEIGHTS => "01",
            SHIFT => 6,
            B => 4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p92_in,
            y(0) => p92_out,
            y(1 to 12 - 1) => dummy92
        );


    p93_in <= x(56) & x(82) & x(202);
    y(93) <= not(p93_out);
    p93 : perceptron
        Generic map (
            WEIGHTS => "000",
            SHIFT => 5,
            B => -9,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p93_in,
            y(0) => p93_out,
            y(1 to 12 - 1) => dummy93
        );


    p94_in(0) <= x(39);
    y(94) <= not(p94_out);
    p94 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => 13,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p94_in,
            y(0) => p94_out,
            y(1 to 12 - 1) => dummy94
        );


    p95_in(0) <= x(249);
    y(95) <= not(p95_out);
    p95 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => -15,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p95_in,
            y(0) => p95_out,
            y(1 to 12 - 1) => dummy95
        );


    p96_in(0) <= x(133);
    y(96) <= not(p96_out);
    p96 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => 11,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p96_in,
            y(0) => p96_out,
            y(1 to 12 - 1) => dummy96
        );


    p97_in <= x(101) & x(116) & x(152);
    y(97) <= not(p97_out);
    p97 : perceptron
        Generic map (
            WEIGHTS => "100",
            SHIFT => 5,
            B => -6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p97_in,
            y(0) => p97_out,
            y(1 to 12 - 1) => dummy97
        );


    p98_in <= x(48) & x(150);
    y(98) <= not(p98_out);
    p98 : perceptron
        Generic map (
            WEIGHTS => "10",
            SHIFT => 6,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p98_in,
            y(0) => p98_out,
            y(1 to 12 - 1) => dummy98
        );


    p99_in <= x(39) & x(133) & x(134) & x(179) & x(213);
    y(99) <= not(p99_out);
    p99 : perceptron
        Generic map (
            WEIGHTS => "00000",
            SHIFT => 6,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p99_in,
            y(0) => p99_out,
            y(1 to 14 - 1) => dummy99
        );


    p100_in <= x(160) & x(213);
    y(100) <= not(p100_out);
    p100 : perceptron
        Generic map (
            WEIGHTS => "00",
            SHIFT => 6,
            B => 7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p100_in,
            y(0) => p100_out,
            y(1 to 12 - 1) => dummy100
        );


    p101_in <= x(65) & x(102) & x(111) & x(150) & x(161) & x(206) & x(244);
    y(101) <= not(p101_out);
    p101 : perceptron
        Generic map (
            WEIGHTS => "1101111",
            SHIFT => 5,
            B => -22,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p101_in,
            y(0) => p101_out,
            y(1 to 13 - 1) => dummy101
        );


    p102_in(0) <= x(63);
    y(102) <= not(p102_out);
    p102 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => 8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p102_in,
            y(0) => p102_out,
            y(1 to 12 - 1) => dummy102
        );


    p103_in <= x(213) & x(239);
    y(103) <= not(p103_out);
    p103 : perceptron
        Generic map (
            WEIGHTS => "10",
            SHIFT => 5,
            B => 12,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p103_in,
            y(0) => p103_out,
            y(1 to 11 - 1) => dummy103
        );


    p104_in <= x(58) & x(69) & x(99) & x(117) & x(150) & x(254);
    y(104) <= not(p104_out);
    p104 : perceptron
        Generic map (
            WEIGHTS => "011001",
            SHIFT => 5,
            B => 7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p104_in,
            y(0) => p104_out,
            y(1 to 13 - 1) => dummy104
        );


    p105_in <= x(150) & x(200) & x(229);
    y(105) <= not(p105_out);
    p105 : perceptron
        Generic map (
            WEIGHTS => "011",
            SHIFT => 6,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p105_in,
            y(0) => p105_out,
            y(1 to 13 - 1) => dummy105
        );


    p106_in <= x(55) & x(222);
    y(106) <= not(p106_out);
    p106 : perceptron
        Generic map (
            WEIGHTS => "10",
            SHIFT => 6,
            B => -7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p106_in,
            y(0) => p106_out,
            y(1 to 12 - 1) => dummy106
        );


    p107_in <= x(104) & x(126) & x(133) & x(150) & x(172) & x(193) & x(200) & x(229) & x(239) & x(246);
    y(107) <= not(p107_out);
    p107 : perceptron
        Generic map (
            WEIGHTS => "0010011100",
            SHIFT => 4,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p107_in,
            y(0) => p107_out,
            y(1 to 13 - 1) => dummy107
        );


    p108_in <= x(101) & x(150);
    y(108) <= not(p108_out);
    p108 : perceptron
        Generic map (
            WEIGHTS => "01",
            SHIFT => 6,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p108_in,
            y(0) => p108_out,
            y(1 to 12 - 1) => dummy108
        );


    p109_in <= x(15) & x(57) & x(69);
    y(109) <= not(p109_out);
    p109 : perceptron
        Generic map (
            WEIGHTS => "000",
            SHIFT => 5,
            B => 4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p109_in,
            y(0) => p109_out,
            y(1 to 12 - 1) => dummy109
        );


    p110_in(0) <= x(150);
    y(110) <= not(p110_out);
    p110 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p110_in,
            y(0) => p110_out,
            y(1 to 12 - 1) => dummy110
        );


    p111_in <= x(12) & x(186);
    y(111) <= not(p111_out);
    p111 : perceptron
        Generic map (
            WEIGHTS => "01",
            SHIFT => 6,
            B => -9,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p111_in,
            y(0) => p111_out,
            y(1 to 12 - 1) => dummy111
        );


    p112_in <= x(93) & x(157) & x(159) & x(177);
    y(112) <= not(p112_out);
    p112 : perceptron
        Generic map (
            WEIGHTS => "1101",
            SHIFT => 6,
            B => 6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p112_in,
            y(0) => p112_out,
            y(1 to 14 - 1) => dummy112
        );


    p113_in(0) <= x(143);
    y(113) <= not(p113_out);
    p113 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p113_in,
            y(0) => p113_out,
            y(1 to 12 - 1) => dummy113
        );


    p114_in <= x(72) & x(229);
    y(114) <= not(p114_out);
    p114 : perceptron
        Generic map (
            WEIGHTS => "10",
            SHIFT => 6,
            B => -20,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p114_in,
            y(0) => p114_out,
            y(1 to 12 - 1) => dummy114
        );


    p115_in <= x(123) & x(175) & x(231) & x(254);
    y(115) <= not(p115_out);
    p115 : perceptron
        Generic map (
            WEIGHTS => "1001",
            SHIFT => 5,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p115_in,
            y(0) => p115_out,
            y(1 to 13 - 1) => dummy115
        );


    p116_in(0) <= x(99);
    y(116) <= not(p116_out);
    p116 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => 22,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p116_in,
            y(0) => p116_out,
            y(1 to 12 - 1) => dummy116
        );


    p117_in(0) <= x(246);
    y(117) <= not(p117_out);
    p117 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => 31,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p117_in,
            y(0) => p117_out,
            y(1 to 12 - 1) => dummy117
        );


    p118_in(0) <= x(95);
    y(118) <= not(p118_out);
    p118 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => -23,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p118_in,
            y(0) => p118_out,
            y(1 to 12 - 1) => dummy118
        );


    p119_in <= x(19) & x(156) & x(163);
    y(119) <= not(p119_out);
    p119 : perceptron
        Generic map (
            WEIGHTS => "000",
            SHIFT => 5,
            B => -34,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p119_in,
            y(0) => p119_out,
            y(1 to 12 - 1) => dummy119
        );


    p120_in(0) <= x(141);
    y(120) <= not(p120_out);
    p120 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 6,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p120_in,
            y(0) => p120_out,
            y(1 to 11 - 1) => dummy120
        );


    p121_in <= x(57) & x(58) & x(74) & x(101) & x(121) & x(133) & x(202) & x(210) & x(241);
    y(121) <= not(p121_out);
    p121 : perceptron
        Generic map (
            WEIGHTS => "100000111",
            SHIFT => 4,
            B => -11,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p121_in,
            y(0) => p121_out,
            y(1 to 13 - 1) => dummy121
        );


    p122_in <= x(99) & x(146) & x(200);
    y(122) <= not(p122_out);
    p122 : perceptron
        Generic map (
            WEIGHTS => "011",
            SHIFT => 5,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p122_in,
            y(0) => p122_out,
            y(1 to 12 - 1) => dummy122
        );


    p123_in <= x(39) & x(85) & x(125);
    y(123) <= not(p123_out);
    p123 : perceptron
        Generic map (
            WEIGHTS => "100",
            SHIFT => 6,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p123_in,
            y(0) => p123_out,
            y(1 to 13 - 1) => dummy123
        );


    p124_in <= x(144) & x(152) & x(176) & x(190) & x(244);
    y(124) <= not(p124_out);
    p124 : perceptron
        Generic map (
            WEIGHTS => "01101",
            SHIFT => 5,
            B => 9,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p124_in,
            y(0) => p124_out,
            y(1 to 13 - 1) => dummy124
        );


    p125_in <= x(78) & x(95) & x(133) & x(215);
    y(125) <= not(p125_out);
    p125 : perceptron
        Generic map (
            WEIGHTS => "0111",
            SHIFT => 5,
            B => -9,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p125_in,
            y(0) => p125_out,
            y(1 to 12 - 1) => dummy125
        );


    p126_in <= x(213) & x(229) & x(239);
    y(126) <= not(p126_out);
    p126 : perceptron
        Generic map (
            WEIGHTS => "110",
            SHIFT => 5,
            B => 9,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p126_in,
            y(0) => p126_out,
            y(1 to 12 - 1) => dummy126
        );


    p127_in <= x(145) & x(244);
    y(127) <= not(p127_out);
    p127 : perceptron
        Generic map (
            WEIGHTS => "00",
            SHIFT => 6,
            B => -20,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p127_in,
            y(0) => p127_out,
            y(1 to 12 - 1) => dummy127
        );


    p128_in <= x(2) & x(89) & x(99) & x(117) & x(150) & x(177) & x(188);
    y(128) <= not(p128_out);
    p128 : perceptron
        Generic map (
            WEIGHTS => "1010000",
            SHIFT => 4,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p128_in,
            y(0) => p128_out,
            y(1 to 12 - 1) => dummy128
        );


    p129_in <= x(37) & x(46) & x(53) & x(63) & x(128) & x(179) & x(233) & x(244);
    y(129) <= not(p129_out);
    p129 : perceptron
        Generic map (
            WEIGHTS => "10110010",
            SHIFT => 5,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p129_in,
            y(0) => p129_out,
            y(1 to 14 - 1) => dummy129
        );


    p130_in <= x(15) & x(99) & x(122) & x(169);
    y(130) <= not(p130_out);
    p130 : perceptron
        Generic map (
            WEIGHTS => "0100",
            SHIFT => 5,
            B => 19,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p130_in,
            y(0) => p130_out,
            y(1 to 12 - 1) => dummy130
        );


    p131_in <= x(40) & x(111) & x(126) & x(172) & x(202);
    y(131) <= not(p131_out);
    p131 : perceptron
        Generic map (
            WEIGHTS => "01000",
            SHIFT => 5,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p131_in,
            y(0) => p131_out,
            y(1 to 13 - 1) => dummy131
        );


    p132_in <= x(101) & x(122) & x(168) & x(188) & x(248);
    y(132) <= not(p132_out);
    p132 : perceptron
        Generic map (
            WEIGHTS => "00001",
            SHIFT => 5,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p132_in,
            y(0) => p132_out,
            y(1 to 13 - 1) => dummy132
        );


    p133_in <= x(25) & x(39);
    y(133) <= not(p133_out);
    p133 : perceptron
        Generic map (
            WEIGHTS => "11",
            SHIFT => 6,
            B => -14,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p133_in,
            y(0) => p133_out,
            y(1 to 12 - 1) => dummy133
        );


    p134_in <= x(14) & x(186);
    y(134) <= not(p134_out);
    p134 : perceptron
        Generic map (
            WEIGHTS => "10",
            SHIFT => 6,
            B => 6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p134_in,
            y(0) => p134_out,
            y(1 to 12 - 1) => dummy134
        );


    p135_in <= x(48) & x(94);
    y(135) <= not(p135_out);
    p135 : perceptron
        Generic map (
            WEIGHTS => "00",
            SHIFT => 6,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p135_in,
            y(0) => p135_out,
            y(1 to 12 - 1) => dummy135
        );


    p136_in(0) <= x(165);
    y(136) <= not(p136_out);
    p136 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p136_in,
            y(0) => p136_out,
            y(1 to 12 - 1) => dummy136
        );


    p137_in <= x(44) & x(111) & x(152) & x(179) & x(244);
    y(137) <= not(p137_out);
    p137 : perceptron
        Generic map (
            WEIGHTS => "11000",
            SHIFT => 5,
            B => -13,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p137_in,
            y(0) => p137_out,
            y(1 to 13 - 1) => dummy137
        );


    p138_in <= x(152) & x(244);
    y(138) <= not(p138_out);
    p138 : perceptron
        Generic map (
            WEIGHTS => "00",
            SHIFT => 6,
            B => -16,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p138_in,
            y(0) => p138_out,
            y(1 to 12 - 1) => dummy138
        );


    p139_in <= x(150) & x(193) & x(200) & x(239);
    y(139) <= not(p139_out);
    p139 : perceptron
        Generic map (
            WEIGHTS => "0110",
            SHIFT => 5,
            B => 6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p139_in,
            y(0) => p139_out,
            y(1 to 13 - 1) => dummy139
        );


    p140_in <= x(101) & x(122) & x(202);
    y(140) <= not(p140_out);
    p140 : perceptron
        Generic map (
            WEIGHTS => "001",
            SHIFT => 6,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p140_in,
            y(0) => p140_out,
            y(1 to 13 - 1) => dummy140
        );


    p141_in <= x(146) & x(156) & x(172) & x(200) & x(239);
    y(141) <= not(p141_out);
    p141 : perceptron
        Generic map (
            WEIGHTS => "01101",
            SHIFT => 5,
            B => -8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p141_in,
            y(0) => p141_out,
            y(1 to 13 - 1) => dummy141
        );


    p142_in(0) <= x(99);
    y(142) <= not(p142_out);
    p142 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => -22,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p142_in,
            y(0) => p142_out,
            y(1 to 12 - 1) => dummy142
        );


    p143_in <= x(90) & x(117) & x(200);
    y(143) <= not(p143_out);
    p143 : perceptron
        Generic map (
            WEIGHTS => "100",
            SHIFT => 5,
            B => -9,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p143_in,
            y(0) => p143_out,
            y(1 to 12 - 1) => dummy143
        );


    p144_in <= x(39) & x(99);
    y(144) <= not(p144_out);
    p144 : perceptron
        Generic map (
            WEIGHTS => "00",
            SHIFT => 7,
            B => -10,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p144_in,
            y(0) => p144_out,
            y(1 to 13 - 1) => dummy144
        );


    p145_in(0) <= x(248);
    y(145) <= not(p145_out);
    p145 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => 4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p145_in,
            y(0) => p145_out,
            y(1 to 12 - 1) => dummy145
        );


    p146_in <= x(116) & x(200);
    y(146) <= not(p146_out);
    p146 : perceptron
        Generic map (
            WEIGHTS => "11",
            SHIFT => 6,
            B => 6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p146_in,
            y(0) => p146_out,
            y(1 to 12 - 1) => dummy146
        );


    p147_in <= x(99) & x(123) & x(156) & x(254);
    y(147) <= not(p147_out);
    p147 : perceptron
        Generic map (
            WEIGHTS => "0000",
            SHIFT => 5,
            B => -23,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p147_in,
            y(0) => p147_out,
            y(1 to 13 - 1) => dummy147
        );


    p148_in <= x(18) & x(63) & x(104) & x(133) & x(134) & x(244);
    y(148) <= not(p148_out);
    p148 : perceptron
        Generic map (
            WEIGHTS => "111000",
            SHIFT => 5,
            B => -14,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p148_in,
            y(0) => p148_out,
            y(1 to 13 - 1) => dummy148
        );


    p149_in(0) <= x(99);
    y(149) <= not(p149_out);
    p149 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => -16,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p149_in,
            y(0) => p149_out,
            y(1 to 12 - 1) => dummy149
        );


    p150_in <= x(63) & x(72) & x(134) & x(144) & x(193);
    y(150) <= not(p150_out);
    p150 : perceptron
        Generic map (
            WEIGHTS => "11011",
            SHIFT => 5,
            B => -10,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p150_in,
            y(0) => p150_out,
            y(1 to 13 - 1) => dummy150
        );


    p151_in <= x(81) & x(172);
    y(151) <= not(p151_out);
    p151 : perceptron
        Generic map (
            WEIGHTS => "00",
            SHIFT => 6,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p151_in,
            y(0) => p151_out,
            y(1 to 12 - 1) => dummy151
        );


    p152_in <= x(116) & x(190);
    y(152) <= not(p152_out);
    p152 : perceptron
        Generic map (
            WEIGHTS => "11",
            SHIFT => 6,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p152_in,
            y(0) => p152_out,
            y(1 to 12 - 1) => dummy152
        );


    p153_in <= x(186) & x(216) & x(243);
    y(153) <= not(p153_out);
    p153 : perceptron
        Generic map (
            WEIGHTS => "100",
            SHIFT => 5,
            B => -12,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p153_in,
            y(0) => p153_out,
            y(1 to 12 - 1) => dummy153
        );


    p154_in <= x(44) & x(122) & x(134) & x(202);
    y(154) <= not(p154_out);
    p154 : perceptron
        Generic map (
            WEIGHTS => "0110",
            SHIFT => 6,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p154_in,
            y(0) => p154_out,
            y(1 to 14 - 1) => dummy154
        );


    p155_in <= x(44) & x(148) & x(186);
    y(155) <= not(p155_out);
    p155 : perceptron
        Generic map (
            WEIGHTS => "111",
            SHIFT => 5,
            B => -8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p155_in,
            y(0) => p155_out,
            y(1 to 12 - 1) => dummy155
        );


    p156_in <= x(51) & x(172);
    y(156) <= not(p156_out);
    p156 : perceptron
        Generic map (
            WEIGHTS => "11",
            SHIFT => 6,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p156_in,
            y(0) => p156_out,
            y(1 to 12 - 1) => dummy156
        );


    p157_in <= x(58) & x(117) & x(188) & x(200) & x(206) & x(224);
    y(157) <= not(p157_out);
    p157 : perceptron
        Generic map (
            WEIGHTS => "111110",
            SHIFT => 5,
            B => -9,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p157_in,
            y(0) => p157_out,
            y(1 to 13 - 1) => dummy157
        );


    p159_in <= x(8) & x(23) & x(108) & x(133) & x(201) & x(224);
    y(159) <= not(p159_out);
    p159 : perceptron
        Generic map (
            WEIGHTS => "101001",
            SHIFT => 4,
            B => -21,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p159_in,
            y(0) => p159_out,
            y(1 to 12 - 1) => dummy159
        );


    p160_in <= x(40) & x(46) & x(81) & x(150) & x(186);
    y(160) <= not(p160_out);
    p160 : perceptron
        Generic map (
            WEIGHTS => "11100",
            SHIFT => 5,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p160_in,
            y(0) => p160_out,
            y(1 to 13 - 1) => dummy160
        );


    p161_in <= x(117) & x(150) & x(243);
    y(161) <= not(p161_out);
    p161 : perceptron
        Generic map (
            WEIGHTS => "001",
            SHIFT => 5,
            B => 6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p161_in,
            y(0) => p161_out,
            y(1 to 12 - 1) => dummy161
        );


    p162_in(0) <= x(3);
    y(162) <= not(p162_out);
    p162 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => -13,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p162_in,
            y(0) => p162_out,
            y(1 to 12 - 1) => dummy162
        );


    p163_in(0) <= x(168);
    y(163) <= not(p163_out);
    p163 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => -15,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p163_in,
            y(0) => p163_out,
            y(1 to 12 - 1) => dummy163
        );


    p164_in <= x(148) & x(186);
    y(164) <= not(p164_out);
    p164 : perceptron
        Generic map (
            WEIGHTS => "00",
            SHIFT => 5,
            B => 8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p164_in,
            y(0) => p164_out,
            y(1 to 11 - 1) => dummy164
        );


    p165_in <= x(19) & x(25);
    y(165) <= not(p165_out);
    p165 : perceptron
        Generic map (
            WEIGHTS => "11",
            SHIFT => 6,
            B => 10,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p165_in,
            y(0) => p165_out,
            y(1 to 12 - 1) => dummy165
        );


    p166_in <= x(144) & x(244);
    y(166) <= not(p166_out);
    p166 : perceptron
        Generic map (
            WEIGHTS => "10",
            SHIFT => 6,
            B => -12,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p166_in,
            y(0) => p166_out,
            y(1 to 12 - 1) => dummy166
        );


    p167_in <= x(5) & x(60) & x(105) & x(116);
    y(167) <= not(p167_out);
    p167 : perceptron
        Generic map (
            WEIGHTS => "1000",
            SHIFT => 5,
            B => -13,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p167_in,
            y(0) => p167_out,
            y(1 to 12 - 1) => dummy167
        );


    p168_in <= x(82) & x(133);
    y(168) <= not(p168_out);
    p168 : perceptron
        Generic map (
            WEIGHTS => "00",
            SHIFT => 6,
            B => -15,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p168_in,
            y(0) => p168_out,
            y(1 to 12 - 1) => dummy168
        );


    p169_in <= x(144) & x(193) & x(244);
    y(169) <= not(p169_out);
    p169 : perceptron
        Generic map (
            WEIGHTS => "100",
            SHIFT => 6,
            B => -10,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p169_in,
            y(0) => p169_out,
            y(1 to 13 - 1) => dummy169
        );


    p170_in <= x(36) & x(177);
    y(170) <= not(p170_out);
    p170 : perceptron
        Generic map (
            WEIGHTS => "11",
            SHIFT => 6,
            B => 4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p170_in,
            y(0) => p170_out,
            y(1 to 12 - 1) => dummy170
        );


    p171_in <= x(44) & x(60) & x(151) & x(193) & x(221);
    y(171) <= not(p171_out);
    p171 : perceptron
        Generic map (
            WEIGHTS => "01010",
            SHIFT => 5,
            B => -9,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p171_in,
            y(0) => p171_out,
            y(1 to 13 - 1) => dummy171
        );


    p172_in <= x(133) & x(193) & x(241);
    y(172) <= not(p172_out);
    p172 : perceptron
        Generic map (
            WEIGHTS => "110",
            SHIFT => 6,
            B => 7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p172_in,
            y(0) => p172_out,
            y(1 to 13 - 1) => dummy172
        );


    p173_in <= x(48) & x(52);
    y(173) <= not(p173_out);
    p173 : perceptron
        Generic map (
            WEIGHTS => "01",
            SHIFT => 6,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p173_in,
            y(0) => p173_out,
            y(1 to 12 - 1) => dummy173
        );


    p174_in <= x(19) & x(67) & x(142) & x(150) & x(188);
    y(174) <= not(p174_out);
    p174 : perceptron
        Generic map (
            WEIGHTS => "00000",
            SHIFT => 5,
            B => -20,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p174_in,
            y(0) => p174_out,
            y(1 to 13 - 1) => dummy174
        );


    p175_in <= x(172) & x(200) & x(229);
    y(175) <= not(p175_out);
    p175 : perceptron
        Generic map (
            WEIGHTS => "100",
            SHIFT => 5,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p175_in,
            y(0) => p175_out,
            y(1 to 12 - 1) => dummy175
        );


    p176_in <= x(44) & x(104) & x(133) & x(150) & x(213) & x(218) & x(244);
    y(176) <= not(p176_out);
    p176 : perceptron
        Generic map (
            WEIGHTS => "0010101",
            SHIFT => 5,
            B => 13,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p176_in,
            y(0) => p176_out,
            y(1 to 13 - 1) => dummy176
        );


    p177_in <= x(48) & x(73) & x(90) & x(98) & x(186) & x(221) & x(235);
    y(177) <= not(p177_out);
    p177 : perceptron
        Generic map (
            WEIGHTS => "0111000",
            SHIFT => 5,
            B => -17,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p177_in,
            y(0) => p177_out,
            y(1 to 13 - 1) => dummy177
        );


    p178_in <= x(62) & x(81) & x(127);
    y(178) <= not(p178_out);
    p178 : perceptron
        Generic map (
            WEIGHTS => "110",
            SHIFT => 6,
            B => -24,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p178_in,
            y(0) => p178_out,
            y(1 to 13 - 1) => dummy178
        );


    p179_in <= x(160) & x(213) & x(222);
    y(179) <= not(p179_out);
    p179 : perceptron
        Generic map (
            WEIGHTS => "001",
            SHIFT => 5,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p179_in,
            y(0) => p179_out,
            y(1 to 12 - 1) => dummy179
        );


    p180_in(0) <= x(39);
    y(180) <= not(p180_out);
    p180 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => 13,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p180_in,
            y(0) => p180_out,
            y(1 to 12 - 1) => dummy180
        );


    p181_in <= x(48) & x(141) & x(159);
    y(181) <= not(p181_out);
    p181 : perceptron
        Generic map (
            WEIGHTS => "011",
            SHIFT => 6,
            B => -8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p181_in,
            y(0) => p181_out,
            y(1 to 13 - 1) => dummy181
        );


    p182_in <= x(21) & x(81) & x(172) & x(182) & x(188) & x(205) & x(215) & x(229) & x(239);
    y(182) <= not(p182_out);
    p182 : perceptron
        Generic map (
            WEIGHTS => "111001001",
            SHIFT => 4,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p182_in,
            y(0) => p182_out,
            y(1 to 13 - 1) => dummy182
        );


    p183_in <= x(97) & x(98) & x(142) & x(177) & x(188);
    y(183) <= not(p183_out);
    p183 : perceptron
        Generic map (
            WEIGHTS => "01000",
            SHIFT => 5,
            B => -11,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p183_in,
            y(0) => p183_out,
            y(1 to 13 - 1) => dummy183
        );


    p184_in <= x(63) & x(82);
    y(184) <= not(p184_out);
    p184 : perceptron
        Generic map (
            WEIGHTS => "00",
            SHIFT => 6,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p184_in,
            y(0) => p184_out,
            y(1 to 12 - 1) => dummy184
        );


    p185_in <= x(104) & x(152) & x(156) & x(172) & x(213) & x(229);
    y(185) <= not(p185_out);
    p185 : perceptron
        Generic map (
            WEIGHTS => "000011",
            SHIFT => 5,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p185_in,
            y(0) => p185_out,
            y(1 to 13 - 1) => dummy185
        );


    p186_in <= x(116) & x(150) & x(152) & x(155) & x(193) & x(198) & x(241) & x(244);
    y(186) <= not(p186_out);
    p186 : perceptron
        Generic map (
            WEIGHTS => "00010010",
            SHIFT => 5,
            B => -22,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p186_in,
            y(0) => p186_out,
            y(1 to 14 - 1) => dummy186
        );


    p187_in <= x(68) & x(228);
    y(187) <= not(p187_out);
    p187 : perceptron
        Generic map (
            WEIGHTS => "01",
            SHIFT => 6,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p187_in,
            y(0) => p187_out,
            y(1 to 12 - 1) => dummy187
        );


    p188_in <= x(111) & x(152) & x(202);
    y(188) <= not(p188_out);
    p188 : perceptron
        Generic map (
            WEIGHTS => "100",
            SHIFT => 6,
            B => -7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p188_in,
            y(0) => p188_out,
            y(1 to 13 - 1) => dummy188
        );


    p189_in <= x(99) & x(172) & x(254);
    y(189) <= not(p189_out);
    p189 : perceptron
        Generic map (
            WEIGHTS => "101",
            SHIFT => 6,
            B => 10,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p189_in,
            y(0) => p189_out,
            y(1 to 13 - 1) => dummy189
        );


    p190_in <= x(26) & x(116) & x(141) & x(220) & x(241) & x(254);
    y(190) <= not(p190_out);
    p190 : perceptron
        Generic map (
            WEIGHTS => "101110",
            SHIFT => 5,
            B => -11,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p190_in,
            y(0) => p190_out,
            y(1 to 13 - 1) => dummy190
        );


    p191_in <= x(40) & x(44) & x(54) & x(114) & x(133) & x(185) & x(190);
    y(191) <= not(p191_out);
    p191 : perceptron
        Generic map (
            WEIGHTS => "0100000",
            SHIFT => 5,
            B => -11,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p191_in,
            y(0) => p191_out,
            y(1 to 13 - 1) => dummy191
        );


    p192_in <= x(74) & x(238);
    y(192) <= not(p192_out);
    p192 : perceptron
        Generic map (
            WEIGHTS => "01",
            SHIFT => 6,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p192_in,
            y(0) => p192_out,
            y(1 to 12 - 1) => dummy192
        );


    p193_in(0) <= x(111);
    y(193) <= not(p193_out);
    p193 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => 8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p193_in,
            y(0) => p193_out,
            y(1 to 12 - 1) => dummy193
        );


    p194_in <= x(60) & x(152);
    y(194) <= not(p194_out);
    p194 : perceptron
        Generic map (
            WEIGHTS => "00",
            SHIFT => 6,
            B => -9,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p194_in,
            y(0) => p194_out,
            y(1 to 12 - 1) => dummy194
        );


    p195_in(0) <= x(39);
    y(195) <= not(p195_out);
    p195 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => 14,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p195_in,
            y(0) => p195_out,
            y(1 to 12 - 1) => dummy195
        );


    p196_in <= x(56) & x(99) & x(134) & x(150) & x(172) & x(177) & x(254);
    y(196) <= not(p196_out);
    p196 : perceptron
        Generic map (
            WEIGHTS => "1110001",
            SHIFT => 5,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p196_in,
            y(0) => p196_out,
            y(1 to 13 - 1) => dummy196
        );


    p197_in <= x(2) & x(56) & x(99) & x(231);
    y(197) <= not(p197_out);
    p197 : perceptron
        Generic map (
            WEIGHTS => "0001",
            SHIFT => 5,
            B => -8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p197_in,
            y(0) => p197_out,
            y(1 to 12 - 1) => dummy197
        );


    p198_in <= x(98) & x(142) & x(150) & x(177) & x(188);
    y(198) <= not(p198_out);
    p198 : perceptron
        Generic map (
            WEIGHTS => "01111",
            SHIFT => 5,
            B => 13,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p198_in,
            y(0) => p198_out,
            y(1 to 13 - 1) => dummy198
        );


    p199_in(0) <= x(200);
    y(199) <= not(p199_out);
    p199 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 6,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p199_in,
            y(0) => p199_out,
            y(1 to 11 - 1) => dummy199
        );


    p200_in <= x(18) & x(152) & x(172) & x(188) & x(193) & x(200) & x(229) & x(239) & x(246);
    y(200) <= not(p200_out);
    p200 : perceptron
        Generic map (
            WEIGHTS => "101000011",
            SHIFT => 5,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p200_in,
            y(0) => p200_out,
            y(1 to 14 - 1) => dummy200
        );


    p201_in <= x(2) & x(45) & x(89) & x(254);
    y(201) <= not(p201_out);
    p201 : perceptron
        Generic map (
            WEIGHTS => "1101",
            SHIFT => 5,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p201_in,
            y(0) => p201_out,
            y(1 to 12 - 1) => dummy201
        );


    p202_in(0) <= x(83);
    y(202) <= not(p202_out);
    p202 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p202_in,
            y(0) => p202_out,
            y(1 to 12 - 1) => dummy202
        );


    p203_in <= x(117) & x(150) & x(186) & x(188);
    y(203) <= not(p203_out);
    p203 : perceptron
        Generic map (
            WEIGHTS => "0000",
            SHIFT => 5,
            B => 6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p203_in,
            y(0) => p203_out,
            y(1 to 13 - 1) => dummy203
        );


    p204_in <= x(77) & x(106) & x(241);
    y(204) <= not(p204_out);
    p204 : perceptron
        Generic map (
            WEIGHTS => "110",
            SHIFT => 6,
            B => 5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p204_in,
            y(0) => p204_out,
            y(1 to 13 - 1) => dummy204
        );


    p205_in <= x(48) & x(97) & x(122);
    y(205) <= not(p205_out);
    p205 : perceptron
        Generic map (
            WEIGHTS => "111",
            SHIFT => 6,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p205_in,
            y(0) => p205_out,
            y(1 to 13 - 1) => dummy205
        );


    p206_in <= x(36) & x(86) & x(169) & x(231);
    y(206) <= not(p206_out);
    p206 : perceptron
        Generic map (
            WEIGHTS => "1000",
            SHIFT => 5,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p206_in,
            y(0) => p206_out,
            y(1 to 12 - 1) => dummy206
        );


    p207_in <= x(40) & x(152) & x(177) & x(186) & x(188);
    y(207) <= not(p207_out);
    p207 : perceptron
        Generic map (
            WEIGHTS => "10000",
            SHIFT => 5,
            B => -13,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p207_in,
            y(0) => p207_out,
            y(1 to 13 - 1) => dummy207
        );


    p208_in <= x(54) & x(78);
    y(208) <= not(p208_out);
    p208 : perceptron
        Generic map (
            WEIGHTS => "10",
            SHIFT => 6,
            B => 8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p208_in,
            y(0) => p208_out,
            y(1 to 12 - 1) => dummy208
        );


    p209_in <= x(44) & x(54) & x(150) & x(193);
    y(209) <= not(p209_out);
    p209 : perceptron
        Generic map (
            WEIGHTS => "0101",
            SHIFT => 5,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p209_in,
            y(0) => p209_out,
            y(1 to 12 - 1) => dummy209
        );


    p210_in <= x(40) & x(119) & x(134) & x(165) & x(179) & x(244);
    y(210) <= not(p210_out);
    p210 : perceptron
        Generic map (
            WEIGHTS => "001011",
            SHIFT => 5,
            B => 7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p210_in,
            y(0) => p210_out,
            y(1 to 13 - 1) => dummy210
        );


    p211_in <= x(39) & x(142) & x(150) & x(188) & x(203);
    y(211) <= not(p211_out);
    p211 : perceptron
        Generic map (
            WEIGHTS => "01110",
            SHIFT => 5,
            B => 18,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p211_in,
            y(0) => p211_out,
            y(1 to 13 - 1) => dummy211
        );


    p212_in <= x(99) & x(129) & x(150) & x(177) & x(250) & x(254);
    y(212) <= not(p212_out);
    p212 : perceptron
        Generic map (
            WEIGHTS => "100001",
            SHIFT => 5,
            B => 7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p212_in,
            y(0) => p212_out,
            y(1 to 13 - 1) => dummy212
        );


    p213_in <= x(89) & x(99) & x(117);
    y(213) <= not(p213_out);
    p213 : perceptron
        Generic map (
            WEIGHTS => "010",
            SHIFT => 5,
            B => 19,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p213_in,
            y(0) => p213_out,
            y(1 to 12 - 1) => dummy213
        );


    p214_in(0) <= x(188);
    y(214) <= not(p214_out);
    p214 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p214_in,
            y(0) => p214_out,
            y(1 to 12 - 1) => dummy214
        );


    p215_in <= x(82) & x(152) & x(244);
    y(215) <= not(p215_out);
    p215 : perceptron
        Generic map (
            WEIGHTS => "100",
            SHIFT => 5,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p215_in,
            y(0) => p215_out,
            y(1 to 12 - 1) => dummy215
        );


    p216_in <= x(12) & x(142) & x(177) & x(188) & x(193) & x(195) & x(200);
    y(216) <= not(p216_out);
    p216 : perceptron
        Generic map (
            WEIGHTS => "0000010",
            SHIFT => 5,
            B => -15,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p216_in,
            y(0) => p216_out,
            y(1 to 13 - 1) => dummy216
        );


    p217_in <= x(36) & x(101) & x(202);
    y(217) <= not(p217_out);
    p217 : perceptron
        Generic map (
            WEIGHTS => "010",
            SHIFT => 6,
            B => 7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p217_in,
            y(0) => p217_out,
            y(1 to 13 - 1) => dummy217
        );


    p218_in <= x(150) & x(193) & x(248);
    y(218) <= not(p218_out);
    p218 : perceptron
        Generic map (
            WEIGHTS => "101",
            SHIFT => 6,
            B => 6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p218_in,
            y(0) => p218_out,
            y(1 to 13 - 1) => dummy218
        );


    p219_in <= x(40) & x(95) & x(133) & x(182);
    y(219) <= not(p219_out);
    p219 : perceptron
        Generic map (
            WEIGHTS => "0000",
            SHIFT => 5,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p219_in,
            y(0) => p219_out,
            y(1 to 12 - 1) => dummy219
        );


    p220_in <= x(81) & x(98) & x(115) & x(142) & x(177) & x(186) & x(188) & x(221);
    y(220) <= not(p220_out);
    p220 : perceptron
        Generic map (
            WEIGHTS => "00011111",
            SHIFT => 4,
            B => 12,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p220_in,
            y(0) => p220_out,
            y(1 to 13 - 1) => dummy220
        );


    p221_in <= x(31) & x(99) & x(254);
    y(221) <= not(p221_out);
    p221 : perceptron
        Generic map (
            WEIGHTS => "000",
            SHIFT => 5,
            B => -11,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p221_in,
            y(0) => p221_out,
            y(1 to 12 - 1) => dummy221
        );


    p222_in <= x(63) & x(244) & x(254);
    y(222) <= not(p222_out);
    p222 : perceptron
        Generic map (
            WEIGHTS => "010",
            SHIFT => 6,
            B => 8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p222_in,
            y(0) => p222_out,
            y(1 to 13 - 1) => dummy222
        );


    p223_in <= x(229) & x(232);
    y(223) <= not(p223_out);
    p223 : perceptron
        Generic map (
            WEIGHTS => "00",
            SHIFT => 6,
            B => -12,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p223_in,
            y(0) => p223_out,
            y(1 to 12 - 1) => dummy223
        );


    p224_in <= x(116) & x(144) & x(152) & x(193) & x(244);
    y(224) <= not(p224_out);
    p224 : perceptron
        Generic map (
            WEIGHTS => "01000",
            SHIFT => 5,
            B => -17,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p224_in,
            y(0) => p224_out,
            y(1 to 13 - 1) => dummy224
        );


    p225_in <= x(39) & x(124);
    y(225) <= not(p225_out);
    p225 : perceptron
        Generic map (
            WEIGHTS => "10",
            SHIFT => 6,
            B => -10,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p225_in,
            y(0) => p225_out,
            y(1 to 12 - 1) => dummy225
        );


    p226_in <= x(39) & x(145) & x(218);
    y(226) <= not(p226_out);
    p226 : perceptron
        Generic map (
            WEIGHTS => "101",
            SHIFT => 6,
            B => -16,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p226_in,
            y(0) => p226_out,
            y(1 to 13 - 1) => dummy226
        );


    p227_in <= x(23) & x(48) & x(120) & x(207);
    y(227) <= not(p227_out);
    p227 : perceptron
        Generic map (
            WEIGHTS => "1001",
            SHIFT => 5,
            B => 13,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p227_in,
            y(0) => p227_out,
            y(1 to 12 - 1) => dummy227
        );


    p228_in <= x(54) & x(129) & x(150);
    y(228) <= not(p228_out);
    p228 : perceptron
        Generic map (
            WEIGHTS => "111",
            SHIFT => 6,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p228_in,
            y(0) => p228_out,
            y(1 to 13 - 1) => dummy228
        );


    p229_in <= x(51) & x(125);
    y(229) <= not(p229_out);
    p229 : perceptron
        Generic map (
            WEIGHTS => "00",
            SHIFT => 6,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p229_in,
            y(0) => p229_out,
            y(1 to 12 - 1) => dummy229
        );


    p230_in <= x(111) & x(131) & x(248);
    y(230) <= not(p230_out);
    p230 : perceptron
        Generic map (
            WEIGHTS => "001",
            SHIFT => 6,
            B => -14,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p230_in,
            y(0) => p230_out,
            y(1 to 13 - 1) => dummy230
        );


    p231_in <= x(44) & x(101);
    y(231) <= not(p231_out);
    p231 : perceptron
        Generic map (
            WEIGHTS => "10",
            SHIFT => 6,
            B => -8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p231_in,
            y(0) => p231_out,
            y(1 to 12 - 1) => dummy231
        );


    p232_in <= x(202) & x(231);
    y(232) <= not(p232_out);
    p232 : perceptron
        Generic map (
            WEIGHTS => "10",
            SHIFT => 5,
            B => 6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p232_in,
            y(0) => p232_out,
            y(1 to 11 - 1) => dummy232
        );


    p233_in <= x(116) & x(194) & x(244);
    y(233) <= not(p233_out);
    p233 : perceptron
        Generic map (
            WEIGHTS => "000",
            SHIFT => 5,
            B => -12,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p233_in,
            y(0) => p233_out,
            y(1 to 12 - 1) => dummy233
        );


    p234_in <= x(39) & x(142) & x(150) & x(221);
    y(234) <= not(p234_out);
    p234 : perceptron
        Generic map (
            WEIGHTS => "1000",
            SHIFT => 5,
            B => -22,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p234_in,
            y(0) => p234_out,
            y(1 to 13 - 1) => dummy234
        );


    p235_in <= x(44) & x(193) & x(224) & x(241);
    y(235) <= not(p235_out);
    p235 : perceptron
        Generic map (
            WEIGHTS => "1011",
            SHIFT => 5,
            B => -12,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p235_in,
            y(0) => p235_out,
            y(1 to 13 - 1) => dummy235
        );


    p236_in <= x(37) & x(106) & x(177);
    y(236) <= not(p236_out);
    p236 : perceptron
        Generic map (
            WEIGHTS => "110",
            SHIFT => 6,
            B => -11,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p236_in,
            y(0) => p236_out,
            y(1 to 13 - 1) => dummy236
        );


    p237_in <= x(90) & x(186) & x(218);
    y(237) <= not(p237_out);
    p237 : perceptron
        Generic map (
            WEIGHTS => "111",
            SHIFT => 5,
            B => -19,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p237_in,
            y(0) => p237_out,
            y(1 to 12 - 1) => dummy237
        );


    p238_in <= x(39) & x(133);
    y(238) <= not(p238_out);
    p238 : perceptron
        Generic map (
            WEIGHTS => "11",
            SHIFT => 6,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p238_in,
            y(0) => p238_out,
            y(1 to 12 - 1) => dummy238
        );


    p239_in(0) <= x(177);
    y(239) <= not(p239_out);
    p239 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => 15,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p239_in,
            y(0) => p239_out,
            y(1 to 12 - 1) => dummy239
        );


    p240_in <= x(172) & x(215);
    y(240) <= not(p240_out);
    p240 : perceptron
        Generic map (
            WEIGHTS => "01",
            SHIFT => 6,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p240_in,
            y(0) => p240_out,
            y(1 to 12 - 1) => dummy240
        );


    p241_in <= x(2) & x(99) & x(117) & x(177) & x(208) & x(228) & x(231) & x(254);
    y(241) <= not(p241_out);
    p241 : perceptron
        Generic map (
            WEIGHTS => "11001101",
            SHIFT => 4,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p241_in,
            y(0) => p241_out,
            y(1 to 13 - 1) => dummy241
        );


    p242_in <= x(111) & x(152) & x(177) & x(188) & x(193) & x(224) & x(239) & x(244);
    y(242) <= not(p242_out);
    p242 : perceptron
        Generic map (
            WEIGHTS => "10000110",
            SHIFT => 5,
            B => -22,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p242_in,
            y(0) => p242_out,
            y(1 to 14 - 1) => dummy242
        );


    p243_in <= x(1) & x(89) & x(117) & x(150) & x(175) & x(254);
    y(243) <= not(p243_out);
    p243 : perceptron
        Generic map (
            WEIGHTS => "100001",
            SHIFT => 4,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p243_in,
            y(0) => p243_out,
            y(1 to 12 - 1) => dummy243
        );


    p244_in <= x(82) & x(94);
    y(244) <= not(p244_out);
    p244 : perceptron
        Generic map (
            WEIGHTS => "00",
            SHIFT => 6,
            B => -11,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p244_in,
            y(0) => p244_out,
            y(1 to 12 - 1) => dummy244
        );


    p245_in <= x(51) & x(54) & x(99) & x(133) & x(172) & x(205);
    y(245) <= not(p245_out);
    p245 : perceptron
        Generic map (
            WEIGHTS => "110011",
            SHIFT => 5,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p245_in,
            y(0) => p245_out,
            y(1 to 13 - 1) => dummy245
        );


    p246_in <= x(60) & x(81);
    y(246) <= not(p246_out);
    p246 : perceptron
        Generic map (
            WEIGHTS => "01",
            SHIFT => 6,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p246_in,
            y(0) => p246_out,
            y(1 to 12 - 1) => dummy246
        );


    p247_in <= x(41) & x(145);
    y(247) <= not(p247_out);
    p247 : perceptron
        Generic map (
            WEIGHTS => "01",
            SHIFT => 5,
            B => 7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p247_in,
            y(0) => p247_out,
            y(1 to 11 - 1) => dummy247
        );


    p248_in <= x(12) & x(23) & x(40) & x(172);
    y(248) <= not(p248_out);
    p248 : perceptron
        Generic map (
            WEIGHTS => "1110",
            SHIFT => 5,
            B => 17,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p248_in,
            y(0) => p248_out,
            y(1 to 12 - 1) => dummy248
        );


    p249_in <= x(148) & x(188) & x(200);
    y(249) <= not(p249_out);
    p249 : perceptron
        Generic map (
            WEIGHTS => "000",
            SHIFT => 6,
            B => 5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p249_in,
            y(0) => p249_out,
            y(1 to 13 - 1) => dummy249
        );


    p250_in <= x(45) & x(94);
    y(250) <= not(p250_out);
    p250 : perceptron
        Generic map (
            WEIGHTS => "00",
            SHIFT => 6,
            B => -14,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p250_in,
            y(0) => p250_out,
            y(1 to 12 - 1) => dummy250
        );


    p251_in <= x(141) & x(160);
    y(251) <= not(p251_out);
    p251 : perceptron
        Generic map (
            WEIGHTS => "00",
            SHIFT => 6,
            B => 8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p251_in,
            y(0) => p251_out,
            y(1 to 12 - 1) => dummy251
        );


    p252_in(0) <= x(126);
    y(252) <= not(p252_out);
    p252 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p252_in,
            y(0) => p252_out,
            y(1 to 12 - 1) => dummy252
        );


    p253_in <= x(24) & x(117) & x(185);
    y(253) <= not(p253_out);
    p253 : perceptron
        Generic map (
            WEIGHTS => "101",
            SHIFT => 5,
            B => 7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p253_in,
            y(0) => p253_out,
            y(1 to 12 - 1) => dummy253
        );


    p254_in <= x(11) & x(99) & x(165) & x(200) & x(222);
    y(254) <= not(p254_out);
    p254 : perceptron
        Generic map (
            WEIGHTS => "10011",
            SHIFT => 5,
            B => 13,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p254_in,
            y(0) => p254_out,
            y(1 to 13 - 1) => dummy254
        );


    p255_in(0) <= x(238);
    y(255) <= not(p255_out);
    p255 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 6,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p255_in,
            y(0) => p255_out,
            y(1 to 11 - 1) => dummy255
        );



end layer_2;

architecture layer_3 of layer is

    Component perceptron
    Generic (
        WEIGHTS : STD_LOGIC_VECTOR := (others => '0');
        SHIFT : Integer;     -- number of shift (left + or right -)
        B : Integer;          -- bias of batch norm
        BATCH_POSITIVE : Boolean    
    );
    Port ( 
        x : in STD_LOGIC_VECTOR;
        y : out STD_LOGIC_VECTOR
   );
    end component;

    -- Signals
    signal p0_in : STD_LOGIC_VECTOR(0 to 7 - 1);
	signal p0_out : STD_LOGIC;
	signal p1_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p1_out : STD_LOGIC;
	signal p2_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p2_out : STD_LOGIC;
	signal p3_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p3_out : STD_LOGIC;
	signal p4_in : STD_LOGIC_VECTOR(0 to 11 - 1);
	signal p4_out : STD_LOGIC;
	signal p5_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p5_out : STD_LOGIC;
	signal p6_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p6_out : STD_LOGIC;
	signal p7_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p7_out : STD_LOGIC;
	signal p8_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p8_out : STD_LOGIC;
	signal p9_in : STD_LOGIC_VECTOR(0 to 7 - 1);
	signal p9_out : STD_LOGIC;
	signal p10_in : STD_LOGIC_VECTOR(0 to 8 - 1);
	signal p10_out : STD_LOGIC;
	signal p11_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p11_out : STD_LOGIC;
	signal p12_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p12_out : STD_LOGIC;
	signal p13_in : STD_LOGIC_VECTOR(0 to 9 - 1);
	signal p13_out : STD_LOGIC;
	signal p14_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p14_out : STD_LOGIC;
	signal p15_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p15_out : STD_LOGIC;
	signal p16_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p16_out : STD_LOGIC;
	signal p17_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p17_out : STD_LOGIC;
	signal p18_in : STD_LOGIC_VECTOR(0 to 7 - 1);
	signal p18_out : STD_LOGIC;
	signal p19_in : STD_LOGIC_VECTOR(0 to 8 - 1);
	signal p19_out : STD_LOGIC;
	signal p20_in : STD_LOGIC_VECTOR(0 to 10 - 1);
	signal p20_out : STD_LOGIC;
	signal p21_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p21_out : STD_LOGIC;
	signal p22_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p22_out : STD_LOGIC;
	signal p23_in : STD_LOGIC_VECTOR(0 to 8 - 1);
	signal p23_out : STD_LOGIC;
	signal p24_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p24_out : STD_LOGIC;
	signal p25_in : STD_LOGIC_VECTOR(0 to 12 - 1);
	signal p25_out : STD_LOGIC;
	signal p26_in : STD_LOGIC_VECTOR(0 to 10 - 1);
	signal p26_out : STD_LOGIC;
	signal p27_in : STD_LOGIC_VECTOR(0 to 8 - 1);
	signal p27_out : STD_LOGIC;
	signal p28_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p28_out : STD_LOGIC;
	signal p29_in : STD_LOGIC_VECTOR(0 to 7 - 1);
	signal p29_out : STD_LOGIC;
	signal p30_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p30_out : STD_LOGIC;
	signal p31_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p31_out : STD_LOGIC;
	signal p32_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p32_out : STD_LOGIC;
	signal p33_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p33_out : STD_LOGIC;
	signal p34_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p34_out : STD_LOGIC;
	signal p35_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p35_out : STD_LOGIC;
	signal p36_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p36_out : STD_LOGIC;
	signal p37_in : STD_LOGIC_VECTOR(0 to 8 - 1);
	signal p37_out : STD_LOGIC;
	signal p38_in : STD_LOGIC_VECTOR(0 to 7 - 1);
	signal p38_out : STD_LOGIC;
	signal p39_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p39_out : STD_LOGIC;
	signal p40_in : STD_LOGIC_VECTOR(0 to 7 - 1);
	signal p40_out : STD_LOGIC;
	signal p41_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p41_out : STD_LOGIC;
	signal p42_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p42_out : STD_LOGIC;
	signal p43_in : STD_LOGIC_VECTOR(0 to 10 - 1);
	signal p43_out : STD_LOGIC;
	signal p44_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p44_out : STD_LOGIC;
	signal p45_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p45_out : STD_LOGIC;
	signal p46_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p46_out : STD_LOGIC;
	signal p47_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p47_out : STD_LOGIC;
	signal p48_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p48_out : STD_LOGIC;
	signal p49_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p49_out : STD_LOGIC;
	signal p50_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p50_out : STD_LOGIC;
	signal p51_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p51_out : STD_LOGIC;
	signal p52_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p52_out : STD_LOGIC;
	signal p53_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p53_out : STD_LOGIC;
	signal p54_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p54_out : STD_LOGIC;
	signal p55_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p55_out : STD_LOGIC;
	signal p56_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p56_out : STD_LOGIC;
	signal p57_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p57_out : STD_LOGIC;
	signal p58_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p58_out : STD_LOGIC;
	signal p59_in : STD_LOGIC_VECTOR(0 to 8 - 1);
	signal p59_out : STD_LOGIC;
	signal p60_in : STD_LOGIC_VECTOR(0 to 12 - 1);
	signal p60_out : STD_LOGIC;
	signal p61_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p61_out : STD_LOGIC;
	signal p62_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p62_out : STD_LOGIC;
	signal p63_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p63_out : STD_LOGIC;
	signal p64_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p64_out : STD_LOGIC;
	signal p65_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p65_out : STD_LOGIC;
	signal p66_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p66_out : STD_LOGIC;
	signal p67_in : STD_LOGIC_VECTOR(0 to 10 - 1);
	signal p67_out : STD_LOGIC;
	signal p68_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p68_out : STD_LOGIC;
	signal p69_in : STD_LOGIC_VECTOR(0 to 9 - 1);
	signal p69_out : STD_LOGIC;
	signal p70_in : STD_LOGIC_VECTOR(0 to 7 - 1);
	signal p70_out : STD_LOGIC;
	signal p71_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p71_out : STD_LOGIC;
	signal p72_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p72_out : STD_LOGIC;
	signal p73_in : STD_LOGIC_VECTOR(0 to 7 - 1);
	signal p73_out : STD_LOGIC;
	signal p74_in : STD_LOGIC_VECTOR(0 to 7 - 1);
	signal p74_out : STD_LOGIC;
	signal p75_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p75_out : STD_LOGIC;
	signal p76_in : STD_LOGIC_VECTOR(0 to 7 - 1);
	signal p76_out : STD_LOGIC;
	signal p77_in : STD_LOGIC_VECTOR(0 to 10 - 1);
	signal p77_out : STD_LOGIC;
	signal p78_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p78_out : STD_LOGIC;
	signal p79_in : STD_LOGIC_VECTOR(0 to 7 - 1);
	signal p79_out : STD_LOGIC;
	signal p80_in : STD_LOGIC_VECTOR(0 to 9 - 1);
	signal p80_out : STD_LOGIC;
	signal p81_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p81_out : STD_LOGIC;
	signal p82_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p82_out : STD_LOGIC;
	signal p83_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p83_out : STD_LOGIC;
	signal p84_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p84_out : STD_LOGIC;
	signal p85_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p85_out : STD_LOGIC;
	signal p86_in : STD_LOGIC_VECTOR(0 to 10 - 1);
	signal p86_out : STD_LOGIC;
	signal p87_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p87_out : STD_LOGIC;
	signal p88_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p88_out : STD_LOGIC;
	signal p89_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p89_out : STD_LOGIC;
	signal p90_in : STD_LOGIC_VECTOR(0 to 8 - 1);
	signal p90_out : STD_LOGIC;
	signal p91_in : STD_LOGIC_VECTOR(0 to 7 - 1);
	signal p91_out : STD_LOGIC;
	signal p92_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p92_out : STD_LOGIC;
	signal p93_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p93_out : STD_LOGIC;
	signal p94_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p94_out : STD_LOGIC;
	signal p95_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p95_out : STD_LOGIC;
	signal p96_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p96_out : STD_LOGIC;
	signal p97_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p97_out : STD_LOGIC;
	signal p98_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p98_out : STD_LOGIC;
	signal p99_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p99_out : STD_LOGIC;
	signal p100_in : STD_LOGIC_VECTOR(0 to 7 - 1);
	signal p100_out : STD_LOGIC;
	signal p101_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p101_out : STD_LOGIC;
	signal p102_in : STD_LOGIC_VECTOR(0 to 12 - 1);
	signal p102_out : STD_LOGIC;
	signal p103_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p103_out : STD_LOGIC;
	signal p104_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p104_out : STD_LOGIC;
	signal p105_in : STD_LOGIC_VECTOR(0 to 8 - 1);
	signal p105_out : STD_LOGIC;
	signal p106_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p106_out : STD_LOGIC;
	signal p107_in : STD_LOGIC_VECTOR(0 to 8 - 1);
	signal p107_out : STD_LOGIC;
	signal p108_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p108_out : STD_LOGIC;
	signal p109_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p109_out : STD_LOGIC;
	signal p110_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p110_out : STD_LOGIC;
	signal p111_in : STD_LOGIC_VECTOR(0 to 7 - 1);
	signal p111_out : STD_LOGIC;
	signal p112_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p112_out : STD_LOGIC;
	signal p113_in : STD_LOGIC_VECTOR(0 to 10 - 1);
	signal p113_out : STD_LOGIC;
	signal p114_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p114_out : STD_LOGIC;
	signal p115_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p115_out : STD_LOGIC;
	signal p116_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p116_out : STD_LOGIC;
	signal p117_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p117_out : STD_LOGIC;
	signal p118_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p118_out : STD_LOGIC;
	signal p119_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p119_out : STD_LOGIC;
	signal p120_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p120_out : STD_LOGIC;
	signal p121_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p121_out : STD_LOGIC;
	signal p122_in : STD_LOGIC_VECTOR(0 to 12 - 1);
	signal p122_out : STD_LOGIC;
	signal p123_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p123_out : STD_LOGIC;
	signal p124_in : STD_LOGIC_VECTOR(0 to 8 - 1);
	signal p124_out : STD_LOGIC;
	signal p125_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p125_out : STD_LOGIC;
	signal p126_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p126_out : STD_LOGIC;
	signal p127_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p127_out : STD_LOGIC;
	signal p128_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p128_out : STD_LOGIC;
	signal p129_in : STD_LOGIC_VECTOR(0 to 8 - 1);
	signal p129_out : STD_LOGIC;
	signal p130_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p130_out : STD_LOGIC;
	signal p131_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p131_out : STD_LOGIC;
	signal p132_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p132_out : STD_LOGIC;
	signal p133_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p133_out : STD_LOGIC;
	signal p134_in : STD_LOGIC_VECTOR(0 to 7 - 1);
	signal p134_out : STD_LOGIC;
	signal p135_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p135_out : STD_LOGIC;
	signal p136_in : STD_LOGIC_VECTOR(0 to 8 - 1);
	signal p136_out : STD_LOGIC;
	signal p137_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p137_out : STD_LOGIC;
	signal p138_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p138_out : STD_LOGIC;
	signal p139_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p139_out : STD_LOGIC;
	signal p140_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p140_out : STD_LOGIC;
	signal p141_in : STD_LOGIC_VECTOR(0 to 8 - 1);
	signal p141_out : STD_LOGIC;
	signal p142_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p142_out : STD_LOGIC;
	signal p143_in : STD_LOGIC_VECTOR(0 to 8 - 1);
	signal p143_out : STD_LOGIC;
	signal p144_in : STD_LOGIC_VECTOR(0 to 7 - 1);
	signal p144_out : STD_LOGIC;
	signal p145_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p145_out : STD_LOGIC;
	signal p146_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p146_out : STD_LOGIC;
	signal p147_in : STD_LOGIC_VECTOR(0 to 8 - 1);
	signal p147_out : STD_LOGIC;
	signal p148_in : STD_LOGIC_VECTOR(0 to 9 - 1);
	signal p148_out : STD_LOGIC;
	signal p149_in : STD_LOGIC_VECTOR(0 to 9 - 1);
	signal p149_out : STD_LOGIC;
	signal p150_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p150_out : STD_LOGIC;
	signal p151_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p151_out : STD_LOGIC;
	signal p152_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p152_out : STD_LOGIC;
	signal p153_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p153_out : STD_LOGIC;
	signal p154_in : STD_LOGIC_VECTOR(0 to 8 - 1);
	signal p154_out : STD_LOGIC;
	signal p155_in : STD_LOGIC_VECTOR(0 to 7 - 1);
	signal p155_out : STD_LOGIC;
	signal p156_in : STD_LOGIC_VECTOR(0 to 7 - 1);
	signal p156_out : STD_LOGIC;
	signal p157_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p157_out : STD_LOGIC;
	signal p158_in : STD_LOGIC_VECTOR(0 to 9 - 1);
	signal p158_out : STD_LOGIC;
	signal p159_in : STD_LOGIC_VECTOR(0 to 9 - 1);
	signal p159_out : STD_LOGIC;
	signal p160_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p160_out : STD_LOGIC;
	signal p161_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p161_out : STD_LOGIC;
	signal p162_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p162_out : STD_LOGIC;
	signal p163_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p163_out : STD_LOGIC;
	signal p164_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p164_out : STD_LOGIC;
	signal p165_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p165_out : STD_LOGIC;
	signal p166_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p166_out : STD_LOGIC;
	signal p167_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p167_out : STD_LOGIC;
	signal p168_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p168_out : STD_LOGIC;
	signal p169_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p169_out : STD_LOGIC;
	signal p170_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p170_out : STD_LOGIC;
	signal p171_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p171_out : STD_LOGIC;
	signal p172_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p172_out : STD_LOGIC;
	signal p173_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p173_out : STD_LOGIC;
	signal p174_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p174_out : STD_LOGIC;
	signal p175_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p175_out : STD_LOGIC;
	signal p176_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p176_out : STD_LOGIC;
	signal p177_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p177_out : STD_LOGIC;
	signal p178_in : STD_LOGIC_VECTOR(0 to 7 - 1);
	signal p178_out : STD_LOGIC;
	signal p179_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p179_out : STD_LOGIC;
	signal p180_in : STD_LOGIC_VECTOR(0 to 10 - 1);
	signal p180_out : STD_LOGIC;
	signal p181_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p181_out : STD_LOGIC;
	signal p182_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p182_out : STD_LOGIC;
	signal p183_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p183_out : STD_LOGIC;
	signal p184_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p184_out : STD_LOGIC;
	signal p185_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p185_out : STD_LOGIC;
	signal p186_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p186_out : STD_LOGIC;
	signal p187_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p187_out : STD_LOGIC;
	signal p188_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p188_out : STD_LOGIC;
	signal p189_in : STD_LOGIC_VECTOR(0 to 10 - 1);
	signal p189_out : STD_LOGIC;
	signal p190_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p190_out : STD_LOGIC;
	signal p191_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p191_out : STD_LOGIC;
	signal p192_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p192_out : STD_LOGIC;
	signal p193_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p193_out : STD_LOGIC;
	signal p194_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p194_out : STD_LOGIC;
	signal p195_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p195_out : STD_LOGIC;
	signal p196_in : STD_LOGIC_VECTOR(0 to 8 - 1);
	signal p196_out : STD_LOGIC;
	signal p197_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p197_out : STD_LOGIC;
	signal p198_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p198_out : STD_LOGIC;
	signal p199_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p199_out : STD_LOGIC;
	signal p200_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p200_out : STD_LOGIC;
	signal p201_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p201_out : STD_LOGIC;
	signal p202_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p202_out : STD_LOGIC;
	signal p203_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p203_out : STD_LOGIC;
	signal p204_in : STD_LOGIC_VECTOR(0 to 7 - 1);
	signal p204_out : STD_LOGIC;
	signal p205_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p205_out : STD_LOGIC;
	signal p206_in : STD_LOGIC_VECTOR(0 to 8 - 1);
	signal p206_out : STD_LOGIC;
	signal p207_in : STD_LOGIC_VECTOR(0 to 7 - 1);
	signal p207_out : STD_LOGIC;
	signal p208_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p208_out : STD_LOGIC;
	signal p209_in : STD_LOGIC_VECTOR(0 to 11 - 1);
	signal p209_out : STD_LOGIC;
	signal p210_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p210_out : STD_LOGIC;
	signal p211_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p211_out : STD_LOGIC;
	signal p212_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p212_out : STD_LOGIC;
	signal p213_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p213_out : STD_LOGIC;
	signal p214_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p214_out : STD_LOGIC;
	signal p215_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p215_out : STD_LOGIC;
	signal p216_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p216_out : STD_LOGIC;
	signal p217_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p217_out : STD_LOGIC;
	signal p218_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p218_out : STD_LOGIC;
	signal p219_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p219_out : STD_LOGIC;
	signal p220_in : STD_LOGIC_VECTOR(0 to 10 - 1);
	signal p220_out : STD_LOGIC;
	signal p222_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p222_out : STD_LOGIC;
	signal p223_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p223_out : STD_LOGIC;
	signal p224_in : STD_LOGIC_VECTOR(0 to 9 - 1);
	signal p224_out : STD_LOGIC;
	signal p225_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p225_out : STD_LOGIC;
	signal p226_in : STD_LOGIC_VECTOR(0 to 10 - 1);
	signal p226_out : STD_LOGIC;
	signal p227_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p227_out : STD_LOGIC;
	signal p228_in : STD_LOGIC_VECTOR(0 to 7 - 1);
	signal p228_out : STD_LOGIC;
	signal p229_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p229_out : STD_LOGIC;
	signal p230_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p230_out : STD_LOGIC;
	signal p231_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p231_out : STD_LOGIC;
	signal p232_in : STD_LOGIC_VECTOR(0 to 8 - 1);
	signal p232_out : STD_LOGIC;
	signal p233_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p233_out : STD_LOGIC;
	signal p234_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p234_out : STD_LOGIC;
	signal p235_in : STD_LOGIC_VECTOR(0 to 8 - 1);
	signal p235_out : STD_LOGIC;
	signal p236_in : STD_LOGIC_VECTOR(0 to 9 - 1);
	signal p236_out : STD_LOGIC;
	signal p237_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p237_out : STD_LOGIC;
	signal p238_in : STD_LOGIC_VECTOR(0 to 9 - 1);
	signal p238_out : STD_LOGIC;
	signal p239_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p239_out : STD_LOGIC;
	signal p240_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p240_out : STD_LOGIC;
	signal p241_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p241_out : STD_LOGIC;
	signal p242_in : STD_LOGIC_VECTOR(0 to 9 - 1);
	signal p242_out : STD_LOGIC;
	signal p243_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p243_out : STD_LOGIC;
	signal p244_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p244_out : STD_LOGIC;
	signal p246_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p246_out : STD_LOGIC;
	signal p247_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p247_out : STD_LOGIC;
	signal p248_in : STD_LOGIC_VECTOR(0 to 9 - 1);
	signal p248_out : STD_LOGIC;
	signal p249_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p249_out : STD_LOGIC;
	signal p250_in : STD_LOGIC_VECTOR(0 to 14 - 1);
	signal p250_out : STD_LOGIC;
	signal p251_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p251_out : STD_LOGIC;
	signal p252_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p252_out : STD_LOGIC;
	signal p253_in : STD_LOGIC_VECTOR(0 to 8 - 1);
	signal p253_out : STD_LOGIC;
	signal p254_in : STD_LOGIC_VECTOR(0 to 9 - 1);
	signal p254_out : STD_LOGIC;
	signal p255_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p255_out : STD_LOGIC;
	
    
    -- Dummies
    signal dummy0 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy1 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy2 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy3 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy4 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy5 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy6 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy7 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy8 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy9 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy10 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy11 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy12 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy13 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy14 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy15 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy16 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy17 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy18 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy19 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy20 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy21 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy22 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy23 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy24 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy25 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy26 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy27 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy28 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy29 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy30 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy31 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy32 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy33 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy34 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy35 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy36 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy37 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy38 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy39 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy40 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy41 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy42 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy43 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy44 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy45 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy46 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy47 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy48 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy49 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy50 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy51 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy52 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy53 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy54 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy55 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy56 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy57 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy58 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy59 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy60 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy61 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy62 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy63 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy64 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy65 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy66 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy67 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy68 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy69 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy70 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy71 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy72 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy73 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy74 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy75 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy76 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy77 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy78 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy79 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy80 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy81 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy82 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy83 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy84 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy85 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy86 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy87 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy88 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy89 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy90 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy91 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy92 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy93 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy94 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy95 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy96 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy97 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy98 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy99 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy100 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy101 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy102 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy103 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy104 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy105 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy106 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy107 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy108 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy109 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy110 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy111 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy112 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy113 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy114 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy115 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy116 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy117 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy118 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy119 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy120 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy121 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy122 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy123 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy124 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy125 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy126 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy127 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy128 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy129 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy130 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy131 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy132 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy133 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy134 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy135 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy136 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy137 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy138 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy139 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy140 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy141 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy142 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy143 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy144 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy145 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy146 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy147 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy148 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy149 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy150 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy151 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy152 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy153 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy154 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy155 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy156 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy157 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy158 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy159 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy160 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy161 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy162 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy163 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy164 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy165 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy166 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy167 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy168 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy169 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy170 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy171 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy172 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy173 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy174 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy175 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy176 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy177 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy178 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy179 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy180 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy181 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy182 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy183 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy184 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy185 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy186 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy187 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy188 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy189 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy190 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy191 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy192 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy193 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy194 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy195 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy196 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy197 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy198 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy199 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy200 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy201 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy202 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy203 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy204 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy205 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy206 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy207 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy208 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy209 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy210 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy211 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy212 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy213 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy214 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy215 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy216 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy217 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy218 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy219 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy220 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy222 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy223 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy224 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy225 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy226 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy227 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy228 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy229 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy230 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy231 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy232 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy233 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy234 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy235 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy236 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy237 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy238 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy239 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy240 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy241 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy242 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy243 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy244 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy246 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy247 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy248 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy249 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy250 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy251 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy252 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy253 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy254 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy255 : STD_LOGIC_VECTOR(0 to 13 - 2);
	 

begin

    
    p0_in <= x(3) & x(66) & x(77) & x(130) & x(174) & x(177) & x(220);
    y(0) <= not(p0_out);
    p0 : perceptron
        Generic map (
            WEIGHTS => "0000001",
            SHIFT => 5,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p0_in,
            y(0) => p0_out,
            y(1 to 13 - 1) => dummy0
        );


    p1_in <= x(43) & x(153) & x(191) & x(194) & x(254);
    y(1) <= not(p1_out);
    p1 : perceptron
        Generic map (
            WEIGHTS => "00001",
            SHIFT => 5,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p1_in,
            y(0) => p1_out,
            y(1 to 13 - 1) => dummy1
        );


    p2_in <= x(153) & x(159) & x(174) & x(229);
    y(2) <= not(p2_out);
    p2 : perceptron
        Generic map (
            WEIGHTS => "1101",
            SHIFT => 6,
            B => 8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p2_in,
            y(0) => p2_out,
            y(1 to 14 - 1) => dummy2
        );


    p3_in <= x(104) & x(170) & x(241);
    y(3) <= not(p3_out);
    p3 : perceptron
        Generic map (
            WEIGHTS => "101",
            SHIFT => 6,
            B => 11,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p3_in,
            y(0) => p3_out,
            y(1 to 13 - 1) => dummy3
        );


    p4_in <= x(5) & x(19) & x(30) & x(43) & x(55) & x(58) & x(159) & x(191) & x(227) & x(235) & x(254);
    y(4) <= not(p4_out);
    p4 : perceptron
        Generic map (
            WEIGHTS => "10000100101",
            SHIFT => 5,
            B => 5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p4_in,
            y(0) => p4_out,
            y(1 to 14 - 1) => dummy4
        );


    p5_in <= x(16) & x(49) & x(50) & x(76) & x(130) & x(170);
    y(5) <= not(p5_out);
    p5 : perceptron
        Generic map (
            WEIGHTS => "110111",
            SHIFT => 5,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p5_in,
            y(0) => p5_out,
            y(1 to 13 - 1) => dummy5
        );


    p6_in <= x(4) & x(14) & x(63) & x(84) & x(101) & x(149);
    y(6) <= not(p6_out);
    p6 : perceptron
        Generic map (
            WEIGHTS => "001001",
            SHIFT => 5,
            B => -11,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p6_in,
            y(0) => p6_out,
            y(1 to 13 - 1) => dummy6
        );


    p7_in <= x(3) & x(34) & x(59);
    y(7) <= not(p7_out);
    p7 : perceptron
        Generic map (
            WEIGHTS => "110",
            SHIFT => 5,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p7_in,
            y(0) => p7_out,
            y(1 to 12 - 1) => dummy7
        );


    p8_in <= x(125) & x(153) & x(191) & x(208) & x(254);
    y(8) <= not(p8_out);
    p8 : perceptron
        Generic map (
            WEIGHTS => "01100",
            SHIFT => 5,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p8_in,
            y(0) => p8_out,
            y(1 to 13 - 1) => dummy8
        );


    p9_in <= x(7) & x(15) & x(76) & x(78) & x(95) & x(230) & x(247);
    y(9) <= not(p9_out);
    p9 : perceptron
        Generic map (
            WEIGHTS => "0110010",
            SHIFT => 5,
            B => 9,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p9_in,
            y(0) => p9_out,
            y(1 to 13 - 1) => dummy9
        );


    p10_in <= x(68) & x(106) & x(114) & x(143) & x(179) & x(190) & x(251) & x(254);
    y(10) <= not(p10_out);
    p10 : perceptron
        Generic map (
            WEIGHTS => "11010100",
            SHIFT => 5,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p10_in,
            y(0) => p10_out,
            y(1 to 14 - 1) => dummy10
        );


    p11_in <= x(143) & x(153) & x(191);
    y(11) <= not(p11_out);
    p11 : perceptron
        Generic map (
            WEIGHTS => "100",
            SHIFT => 6,
            B => 10,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p11_in,
            y(0) => p11_out,
            y(1 to 13 - 1) => dummy11
        );


    p12_in <= x(22) & x(66) & x(98) & x(114) & x(179) & x(227);
    y(12) <= not(p12_out);
    p12 : perceptron
        Generic map (
            WEIGHTS => "110001",
            SHIFT => 5,
            B => -7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p12_in,
            y(0) => p12_out,
            y(1 to 13 - 1) => dummy12
        );


    p13_in <= x(16) & x(50) & x(91) & x(159) & x(191) & x(205) & x(227) & x(231) & x(248);
    y(13) <= not(p13_out);
    p13 : perceptron
        Generic map (
            WEIGHTS => "011111010",
            SHIFT => 4,
            B => 4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p13_in,
            y(0) => p13_out,
            y(1 to 13 - 1) => dummy13
        );


    p14_in <= x(109) & x(125) & x(128) & x(159) & x(191);
    y(14) <= not(p14_out);
    p14 : perceptron
        Generic map (
            WEIGHTS => "00111",
            SHIFT => 5,
            B => -6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p14_in,
            y(0) => p14_out,
            y(1 to 13 - 1) => dummy14
        );


    p15_in <= x(116) & x(125) & x(191) & x(208) & x(232) & x(254);
    y(15) <= not(p15_out);
    p15 : perceptron
        Generic map (
            WEIGHTS => "010101",
            SHIFT => 5,
            B => -11,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p15_in,
            y(0) => p15_out,
            y(1 to 13 - 1) => dummy15
        );


    p16_in <= x(121) & x(125) & x(164) & x(237);
    y(16) <= not(p16_out);
    p16 : perceptron
        Generic map (
            WEIGHTS => "1001",
            SHIFT => 5,
            B => -6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p16_in,
            y(0) => p16_out,
            y(1 to 13 - 1) => dummy16
        );


    p17_in <= x(43) & x(191) & x(254);
    y(17) <= not(p17_out);
    p17 : perceptron
        Generic map (
            WEIGHTS => "110",
            SHIFT => 6,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p17_in,
            y(0) => p17_out,
            y(1 to 13 - 1) => dummy17
        );


    p18_in <= x(3) & x(66) & x(77) & x(121) & x(190) & x(232) & x(254);
    y(18) <= not(p18_out);
    p18 : perceptron
        Generic map (
            WEIGHTS => "1111011",
            SHIFT => 5,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p18_in,
            y(0) => p18_out,
            y(1 to 13 - 1) => dummy18
        );


    p19_in <= x(13) & x(15) & x(61) & x(77) & x(79) & x(177) & x(191) & x(204);
    y(19) <= not(p19_out);
    p19 : perceptron
        Generic map (
            WEIGHTS => "01000010",
            SHIFT => 5,
            B => -8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p19_in,
            y(0) => p19_out,
            y(1 to 14 - 1) => dummy19
        );


    p20_in <= x(3) & x(13) & x(30) & x(37) & x(59) & x(66) & x(155) & x(164) & x(214) & x(255);
    y(20) <= not(p20_out);
    p20 : perceptron
        Generic map (
            WEIGHTS => "0011100100",
            SHIFT => 4,
            B => 5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p20_in,
            y(0) => p20_out,
            y(1 to 13 - 1) => dummy20
        );


    p21_in <= x(5) & x(43) & x(96) & x(227) & x(239) & x(254);
    y(21) <= not(p21_out);
    p21 : perceptron
        Generic map (
            WEIGHTS => "010000",
            SHIFT => 5,
            B => -8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p21_in,
            y(0) => p21_out,
            y(1 to 13 - 1) => dummy21
        );


    p22_in <= x(93) & x(153) & x(191) & x(208) & x(241) & x(243);
    y(22) <= not(p22_out);
    p22 : perceptron
        Generic map (
            WEIGHTS => "111000",
            SHIFT => 5,
            B => -7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p22_in,
            y(0) => p22_out,
            y(1 to 13 - 1) => dummy22
        );


    p23_in <= x(32) & x(43) & x(77) & x(101) & x(104) & x(248) & x(253) & x(254);
    y(23) <= not(p23_out);
    p23 : perceptron
        Generic map (
            WEIGHTS => "11110000",
            SHIFT => 5,
            B => 12,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p23_in,
            y(0) => p23_out,
            y(1 to 14 - 1) => dummy23
        );


    p24_in(0) <= x(191);
    y(24) <= not(p24_out);
    p24 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => -9,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p24_in,
            y(0) => p24_out,
            y(1 to 12 - 1) => dummy24
        );


    p25_in <= x(3) & x(34) & x(43) & x(68) & x(115) & x(121) & x(143) & x(146) & x(157) & x(159) & x(241) & x(248);
    y(25) <= not(p25_out);
    p25 : perceptron
        Generic map (
            WEIGHTS => "010000011001",
            SHIFT => 4,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p25_in,
            y(0) => p25_out,
            y(1 to 13 - 1) => dummy25
        );


    p26_in <= x(13) & x(37) & x(62) & x(112) & x(115) & x(127) & x(134) & x(190) & x(237) & x(241);
    y(26) <= not(p26_out);
    p26 : perceptron
        Generic map (
            WEIGHTS => "0010011100",
            SHIFT => 5,
            B => 4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p26_in,
            y(0) => p26_out,
            y(1 to 14 - 1) => dummy26
        );


    p27_in <= x(41) & x(131) & x(170) & x(208) & x(220) & x(228) & x(236) & x(241);
    y(27) <= not(p27_out);
    p27 : perceptron
        Generic map (
            WEIGHTS => "11001011",
            SHIFT => 5,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p27_in,
            y(0) => p27_out,
            y(1 to 14 - 1) => dummy27
        );


    p28_in <= x(77) & x(193) & x(232);
    y(28) <= not(p28_out);
    p28 : perceptron
        Generic map (
            WEIGHTS => "101",
            SHIFT => 6,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p28_in,
            y(0) => p28_out,
            y(1 to 13 - 1) => dummy28
        );


    p29_in <= x(3) & x(90) & x(109) & x(153) & x(187) & x(235) & x(255);
    y(29) <= not(p29_out);
    p29 : perceptron
        Generic map (
            WEIGHTS => "0111101",
            SHIFT => 5,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p29_in,
            y(0) => p29_out,
            y(1 to 13 - 1) => dummy29
        );


    p30_in <= x(87) & x(101) & x(202) & x(230) & x(231);
    y(30) <= not(p30_out);
    p30 : perceptron
        Generic map (
            WEIGHTS => "01110",
            SHIFT => 5,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p30_in,
            y(0) => p30_out,
            y(1 to 13 - 1) => dummy30
        );


    p31_in <= x(8) & x(118) & x(254);
    y(31) <= not(p31_out);
    p31 : perceptron
        Generic map (
            WEIGHTS => "010",
            SHIFT => 5,
            B => -10,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p31_in,
            y(0) => p31_out,
            y(1 to 12 - 1) => dummy31
        );


    p32_in <= x(19) & x(101) & x(113) & x(170) & x(208) & x(253);
    y(32) <= not(p32_out);
    p32 : perceptron
        Generic map (
            WEIGHTS => "111000",
            SHIFT => 5,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p32_in,
            y(0) => p32_out,
            y(1 to 13 - 1) => dummy32
        );


    p33_in <= x(16) & x(66) & x(68) & x(232);
    y(33) <= not(p33_out);
    p33 : perceptron
        Generic map (
            WEIGHTS => "0010",
            SHIFT => 5,
            B => -6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p33_in,
            y(0) => p33_out,
            y(1 to 12 - 1) => dummy33
        );


    p34_in <= x(43) & x(77) & x(205) & x(208) & x(241);
    y(34) <= not(p34_out);
    p34 : perceptron
        Generic map (
            WEIGHTS => "00110",
            SHIFT => 5,
            B => -17,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p34_in,
            y(0) => p34_out,
            y(1 to 13 - 1) => dummy34
        );


    p35_in <= x(43) & x(59) & x(135) & x(190) & x(241) & x(254);
    y(35) <= not(p35_out);
    p35 : perceptron
        Generic map (
            WEIGHTS => "111110",
            SHIFT => 5,
            B => 6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p35_in,
            y(0) => p35_out,
            y(1 to 13 - 1) => dummy35
        );


    p36_in <= x(61) & x(79) & x(114) & x(190) & x(251) & x(254);
    y(36) <= not(p36_out);
    p36 : perceptron
        Generic map (
            WEIGHTS => "110100",
            SHIFT => 5,
            B => 5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p36_in,
            y(0) => p36_out,
            y(1 to 13 - 1) => dummy36
        );


    p37_in <= x(8) & x(15) & x(63) & x(115) & x(119) & x(229) & x(241) & x(254);
    y(37) <= not(p37_out);
    p37 : perceptron
        Generic map (
            WEIGHTS => "11010110",
            SHIFT => 5,
            B => 17,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p37_in,
            y(0) => p37_out,
            y(1 to 14 - 1) => dummy37
        );


    p38_in <= x(3) & x(13) & x(89) & x(159) & x(177) & x(191) & x(205);
    y(38) <= not(p38_out);
    p38 : perceptron
        Generic map (
            WEIGHTS => "1110100",
            SHIFT => 5,
            B => 5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p38_in,
            y(0) => p38_out,
            y(1 to 13 - 1) => dummy38
        );


    p39_in <= x(33) & x(106) & x(136) & x(232);
    y(39) <= not(p39_out);
    p39 : perceptron
        Generic map (
            WEIGHTS => "1000",
            SHIFT => 5,
            B => -11,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p39_in,
            y(0) => p39_out,
            y(1 to 13 - 1) => dummy39
        );


    p40_in <= x(70) & x(86) & x(101) & x(149) & x(202) & x(228) & x(229);
    y(40) <= not(p40_out);
    p40 : perceptron
        Generic map (
            WEIGHTS => "1010101",
            SHIFT => 4,
            B => 13,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p40_in,
            y(0) => p40_out,
            y(1 to 12 - 1) => dummy40
        );


    p41_in <= x(3) & x(43) & x(77) & x(90) & x(177) & x(241);
    y(41) <= not(p41_out);
    p41 : perceptron
        Generic map (
            WEIGHTS => "111011",
            SHIFT => 5,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p41_in,
            y(0) => p41_out,
            y(1 to 13 - 1) => dummy41
        );


    p42_in <= x(102) & x(105) & x(127) & x(154) & x(191);
    y(42) <= not(p42_out);
    p42 : perceptron
        Generic map (
            WEIGHTS => "10010",
            SHIFT => 5,
            B => -11,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p42_in,
            y(0) => p42_out,
            y(1 to 13 - 1) => dummy42
        );


    p43_in <= x(22) & x(106) & x(114) & x(120) & x(135) & x(167) & x(190) & x(233) & x(251) & x(254);
    y(43) <= not(p43_out);
    p43 : perceptron
        Generic map (
            WEIGHTS => "0010000011",
            SHIFT => 4,
            B => -13,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p43_in,
            y(0) => p43_out,
            y(1 to 13 - 1) => dummy43
        );


    p44_in <= x(30) & x(155) & x(164) & x(248);
    y(44) <= not(p44_out);
    p44 : perceptron
        Generic map (
            WEIGHTS => "0100",
            SHIFT => 5,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p44_in,
            y(0) => p44_out,
            y(1 to 13 - 1) => dummy44
        );


    p45_in <= x(13) & x(18) & x(66) & x(68) & x(146) & x(159);
    y(45) <= not(p45_out);
    p45 : perceptron
        Generic map (
            WEIGHTS => "101010",
            SHIFT => 5,
            B => 8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p45_in,
            y(0) => p45_out,
            y(1 to 13 - 1) => dummy45
        );


    p46_in <= x(178) & x(232) & x(241);
    y(46) <= not(p46_out);
    p46 : perceptron
        Generic map (
            WEIGHTS => "000",
            SHIFT => 6,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p46_in,
            y(0) => p46_out,
            y(1 to 13 - 1) => dummy46
        );


    p47_in <= x(112) & x(115) & x(127) & x(155) & x(191) & x(241);
    y(47) <= not(p47_out);
    p47 : perceptron
        Generic map (
            WEIGHTS => "110101",
            SHIFT => 5,
            B => -13,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p47_in,
            y(0) => p47_out,
            y(1 to 13 - 1) => dummy47
        );


    p48_in <= x(41) & x(101) & x(149) & x(230);
    y(48) <= not(p48_out);
    p48 : perceptron
        Generic map (
            WEIGHTS => "1101",
            SHIFT => 5,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p48_in,
            y(0) => p48_out,
            y(1 to 13 - 1) => dummy48
        );


    p49_in <= x(3) & x(30) & x(194) & x(255);
    y(49) <= not(p49_out);
    p49 : perceptron
        Generic map (
            WEIGHTS => "0110",
            SHIFT => 6,
            B => 11,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p49_in,
            y(0) => p49_out,
            y(1 to 13 - 1) => dummy49
        );


    p50_in <= x(118) & x(187) & x(203);
    y(50) <= not(p50_out);
    p50 : perceptron
        Generic map (
            WEIGHTS => "001",
            SHIFT => 6,
            B => 8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p50_in,
            y(0) => p50_out,
            y(1 to 13 - 1) => dummy50
        );


    p51_in <= x(41) & x(115) & x(121) & x(125) & x(208) & x(241);
    y(51) <= not(p51_out);
    p51 : perceptron
        Generic map (
            WEIGHTS => "111001",
            SHIFT => 5,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p51_in,
            y(0) => p51_out,
            y(1 to 13 - 1) => dummy51
        );


    p52_in <= x(49) & x(74) & x(76) & x(81) & x(131) & x(232);
    y(52) <= not(p52_out);
    p52 : perceptron
        Generic map (
            WEIGHTS => "000010",
            SHIFT => 5,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p52_in,
            y(0) => p52_out,
            y(1 to 13 - 1) => dummy52
        );


    p53_in <= x(87) & x(101) & x(104) & x(109) & x(164) & x(244);
    y(53) <= not(p53_out);
    p53 : perceptron
        Generic map (
            WEIGHTS => "101000",
            SHIFT => 5,
            B => -13,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p53_in,
            y(0) => p53_out,
            y(1 to 13 - 1) => dummy53
        );


    p54_in <= x(104) & x(190) & x(237);
    y(54) <= not(p54_out);
    p54 : perceptron
        Generic map (
            WEIGHTS => "101",
            SHIFT => 6,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p54_in,
            y(0) => p54_out,
            y(1 to 13 - 1) => dummy54
        );


    p55_in <= x(153) & x(237);
    y(55) <= not(p55_out);
    p55 : perceptron
        Generic map (
            WEIGHTS => "10",
            SHIFT => 7,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p55_in,
            y(0) => p55_out,
            y(1 to 13 - 1) => dummy55
        );


    p56_in <= x(22) & x(48) & x(106) & x(114) & x(188) & x(251);
    y(56) <= not(p56_out);
    p56 : perceptron
        Generic map (
            WEIGHTS => "000101",
            SHIFT => 5,
            B => -12,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p56_in,
            y(0) => p56_out,
            y(1 to 13 - 1) => dummy56
        );


    p57_in <= x(15) & x(87) & x(222);
    y(57) <= not(p57_out);
    p57 : perceptron
        Generic map (
            WEIGHTS => "101",
            SHIFT => 6,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p57_in,
            y(0) => p57_out,
            y(1 to 13 - 1) => dummy57
        );


    p58_in <= x(32) & x(43) & x(104) & x(232) & x(248) & x(254);
    y(58) <= not(p58_out);
    p58 : perceptron
        Generic map (
            WEIGHTS => "001011",
            SHIFT => 5,
            B => -12,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p58_in,
            y(0) => p58_out,
            y(1 to 13 - 1) => dummy58
        );


    p59_in <= x(8) & x(13) & x(159) & x(184) & x(191) & x(227) & x(235) & x(248);
    y(59) <= not(p59_out);
    p59 : perceptron
        Generic map (
            WEIGHTS => "10111010",
            SHIFT => 4,
            B => 6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p59_in,
            y(0) => p59_out,
            y(1 to 13 - 1) => dummy59
        );


    p60_in <= x(10) & x(41) & x(59) & x(61) & x(71) & x(89) & x(92) & x(98) & x(129) & x(152) & x(190) & x(241);
    y(60) <= not(p60_out);
    p60 : perceptron
        Generic map (
            WEIGHTS => "101111000010",
            SHIFT => 5,
            B => 4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p60_in,
            y(0) => p60_out,
            y(1 to 14 - 1) => dummy60
        );


    p61_in <= x(66) & x(109) & x(123) & x(178);
    y(61) <= not(p61_out);
    p61 : perceptron
        Generic map (
            WEIGHTS => "1110",
            SHIFT => 6,
            B => 8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p61_in,
            y(0) => p61_out,
            y(1 to 14 - 1) => dummy61
        );


    p62_in <= x(3) & x(36) & x(164) & x(232);
    y(62) <= not(p62_out);
    p62 : perceptron
        Generic map (
            WEIGHTS => "0110",
            SHIFT => 5,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p62_in,
            y(0) => p62_out,
            y(1 to 12 - 1) => dummy62
        );


    p63_in <= x(208) & x(243);
    y(63) <= not(p63_out);
    p63 : perceptron
        Generic map (
            WEIGHTS => "00",
            SHIFT => 6,
            B => 13,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p63_in,
            y(0) => p63_out,
            y(1 to 12 - 1) => dummy63
        );


    p64_in <= x(49) & x(232);
    y(64) <= not(p64_out);
    p64 : perceptron
        Generic map (
            WEIGHTS => "00",
            SHIFT => 6,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p64_in,
            y(0) => p64_out,
            y(1 to 12 - 1) => dummy64
        );


    p65_in <= x(52) & x(87) & x(202) & x(230) & x(255);
    y(65) <= not(p65_out);
    p65 : perceptron
        Generic map (
            WEIGHTS => "01000",
            SHIFT => 5,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p65_in,
            y(0) => p65_out,
            y(1 to 13 - 1) => dummy65
        );


    p66_in <= x(47) & x(49) & x(74) & x(81) & x(131) & x(232);
    y(66) <= not(p66_out);
    p66 : perceptron
        Generic map (
            WEIGHTS => "111101",
            SHIFT => 5,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p66_in,
            y(0) => p66_out,
            y(1 to 13 - 1) => dummy66
        );


    p67_in <= x(13) & x(34) & x(125) & x(141) & x(159) & x(172) & x(191) & x(227) & x(241) & x(248);
    y(67) <= not(p67_out);
    p67 : perceptron
        Generic map (
            WEIGHTS => "0001101000",
            SHIFT => 4,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p67_in,
            y(0) => p67_out,
            y(1 to 13 - 1) => dummy67
        );


    p68_in <= x(101) & x(104) & x(229) & x(246) & x(253);
    y(68) <= not(p68_out);
    p68 : perceptron
        Generic map (
            WEIGHTS => "01111",
            SHIFT => 5,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p68_in,
            y(0) => p68_out,
            y(1 to 13 - 1) => dummy68
        );


    p69_in <= x(26) & x(34) & x(43) & x(68) & x(104) & x(159) & x(191) & x(235) & x(254);
    y(69) <= not(p69_out);
    p69 : perceptron
        Generic map (
            WEIGHTS => "101101110",
            SHIFT => 5,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p69_in,
            y(0) => p69_out,
            y(1 to 14 - 1) => dummy69
        );


    p70_in <= x(41) & x(104) & x(115) & x(121) & x(125) & x(241) & x(243);
    y(70) <= not(p70_out);
    p70 : perceptron
        Generic map (
            WEIGHTS => "1111011",
            SHIFT => 5,
            B => -7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p70_in,
            y(0) => p70_out,
            y(1 to 13 - 1) => dummy70
        );


    p71_in <= x(30) & x(43) & x(66) & x(131);
    y(71) <= not(p71_out);
    p71 : perceptron
        Generic map (
            WEIGHTS => "0011",
            SHIFT => 5,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p71_in,
            y(0) => p71_out,
            y(1 to 12 - 1) => dummy71
        );


    p72_in <= x(194) & x(248);
    y(72) <= not(p72_out);
    p72 : perceptron
        Generic map (
            WEIGHTS => "00",
            SHIFT => 6,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p72_in,
            y(0) => p72_out,
            y(1 to 12 - 1) => dummy72
        );


    p73_in <= x(30) & x(37) & x(44) & x(94) & x(101) & x(229) & x(235);
    y(73) <= not(p73_out);
    p73 : perceptron
        Generic map (
            WEIGHTS => "1001011",
            SHIFT => 5,
            B => 13,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p73_in,
            y(0) => p73_out,
            y(1 to 13 - 1) => dummy73
        );


    p74_in <= x(13) & x(66) & x(68) & x(141) & x(159) & x(227) & x(248);
    y(74) <= not(p74_out);
    p74 : perceptron
        Generic map (
            WEIGHTS => "1100011",
            SHIFT => 5,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p74_in,
            y(0) => p74_out,
            y(1 to 13 - 1) => dummy74
        );


    p75_in <= x(30) & x(153) & x(208);
    y(75) <= not(p75_out);
    p75 : perceptron
        Generic map (
            WEIGHTS => "101",
            SHIFT => 5,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p75_in,
            y(0) => p75_out,
            y(1 to 12 - 1) => dummy75
        );


    p76_in <= x(125) & x(153) & x(155) & x(191) & x(199) & x(208) & x(215);
    y(76) <= not(p76_out);
    p76 : perceptron
        Generic map (
            WEIGHTS => "0111101",
            SHIFT => 5,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p76_in,
            y(0) => p76_out,
            y(1 to 13 - 1) => dummy76
        );


    p77_in <= x(3) & x(13) & x(14) & x(77) & x(85) & x(90) & x(160) & x(174) & x(237) & x(248);
    y(77) <= not(p77_out);
    p77 : perceptron
        Generic map (
            WEIGHTS => "1111001101",
            SHIFT => 5,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p77_in,
            y(0) => p77_out,
            y(1 to 14 - 1) => dummy77
        );


    p78_in <= x(188) & x(191) & x(206) & x(232);
    y(78) <= not(p78_out);
    p78 : perceptron
        Generic map (
            WEIGHTS => "1000",
            SHIFT => 5,
            B => 5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p78_in,
            y(0) => p78_out,
            y(1 to 13 - 1) => dummy78
        );


    p79_in <= x(8) & x(82) & x(124) & x(129) & x(229) & x(241) & x(254);
    y(79) <= not(p79_out);
    p79 : perceptron
        Generic map (
            WEIGHTS => "1010001",
            SHIFT => 5,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p79_in,
            y(0) => p79_out,
            y(1 to 13 - 1) => dummy79
        );


    p80_in <= x(43) & x(59) & x(118) & x(121) & x(125) & x(155) & x(164) & x(199) & x(237);
    y(80) <= not(p80_out);
    p80 : perceptron
        Generic map (
            WEIGHTS => "111010100",
            SHIFT => 4,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p80_in,
            y(0) => p80_out,
            y(1 to 13 - 1) => dummy80
        );


    p81_in <= x(3) & x(49) & x(101) & x(174) & x(220) & x(248);
    y(81) <= not(p81_out);
    p81 : perceptron
        Generic map (
            WEIGHTS => "110101",
            SHIFT => 5,
            B => -14,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p81_in,
            y(0) => p81_out,
            y(1 to 13 - 1) => dummy81
        );


    p82_in <= x(179) & x(246);
    y(82) <= not(p82_out);
    p82 : perceptron
        Generic map (
            WEIGHTS => "00",
            SHIFT => 6,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p82_in,
            y(0) => p82_out,
            y(1 to 12 - 1) => dummy82
        );


    p83_in <= x(13) & x(29) & x(131) & x(190) & x(241) & x(254);
    y(83) <= not(p83_out);
    p83 : perceptron
        Generic map (
            WEIGHTS => "100011",
            SHIFT => 5,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p83_in,
            y(0) => p83_out,
            y(1 to 13 - 1) => dummy83
        );


    p84_in <= x(28) & x(90) & x(101) & x(153) & x(157) & x(246);
    y(84) <= not(p84_out);
    p84 : perceptron
        Generic map (
            WEIGHTS => "011110",
            SHIFT => 5,
            B => -6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p84_in,
            y(0) => p84_out,
            y(1 to 13 - 1) => dummy84
        );


    p85_in <= x(104) & x(118) & x(125) & x(191) & x(215) & x(240);
    y(85) <= not(p85_out);
    p85 : perceptron
        Generic map (
            WEIGHTS => "100100",
            SHIFT => 5,
            B => 6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p85_in,
            y(0) => p85_out,
            y(1 to 13 - 1) => dummy85
        );


    p86_in <= x(3) & x(25) & x(43) & x(77) & x(117) & x(151) & x(159) & x(177) & x(240) & x(254);
    y(86) <= not(p86_out);
    p86 : perceptron
        Generic map (
            WEIGHTS => "0100010011",
            SHIFT => 5,
            B => -13,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p86_in,
            y(0) => p86_out,
            y(1 to 14 - 1) => dummy86
        );


    p87_in <= x(101) & x(215);
    y(87) <= not(p87_out);
    p87 : perceptron
        Generic map (
            WEIGHTS => "00",
            SHIFT => 6,
            B => 5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p87_in,
            y(0) => p87_out,
            y(1 to 12 - 1) => dummy87
        );


    p88_in <= x(43) & x(113) & x(115) & x(157) & x(241);
    y(88) <= not(p88_out);
    p88 : perceptron
        Generic map (
            WEIGHTS => "11101",
            SHIFT => 5,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p88_in,
            y(0) => p88_out,
            y(1 to 13 - 1) => dummy88
        );


    p89_in <= x(153) & x(208);
    y(89) <= not(p89_out);
    p89 : perceptron
        Generic map (
            WEIGHTS => "01",
            SHIFT => 6,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p89_in,
            y(0) => p89_out,
            y(1 to 12 - 1) => dummy89
        );


    p90_in <= x(13) & x(26) & x(104) & x(115) & x(229) & x(237) & x(241) & x(243);
    y(90) <= not(p90_out);
    p90 : perceptron
        Generic map (
            WEIGHTS => "10111111",
            SHIFT => 4,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p90_in,
            y(0) => p90_out,
            y(1 to 13 - 1) => dummy90
        );


    p91_in <= x(18) & x(66) & x(68) & x(128) & x(143) & x(153) & x(208);
    y(91) <= not(p91_out);
    p91 : perceptron
        Generic map (
            WEIGHTS => "1011101",
            SHIFT => 5,
            B => -7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p91_in,
            y(0) => p91_out,
            y(1 to 13 - 1) => dummy91
        );


    p92_in <= x(43) & x(241);
    y(92) <= not(p92_out);
    p92 : perceptron
        Generic map (
            WEIGHTS => "11",
            SHIFT => 6,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p92_in,
            y(0) => p92_out,
            y(1 to 12 - 1) => dummy92
        );


    p93_in <= x(3) & x(30) & x(43) & x(177) & x(220) & x(246);
    y(93) <= not(p93_out);
    p93 : perceptron
        Generic map (
            WEIGHTS => "000010",
            SHIFT => 5,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p93_in,
            y(0) => p93_out,
            y(1 to 13 - 1) => dummy93
        );


    p94_in <= x(1) & x(22) & x(164) & x(165) & x(248);
    y(94) <= not(p94_out);
    p94 : perceptron
        Generic map (
            WEIGHTS => "00010",
            SHIFT => 5,
            B => -13,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p94_in,
            y(0) => p94_out,
            y(1 to 13 - 1) => dummy94
        );


    p95_in <= x(6) & x(41) & x(160) & x(235) & x(237);
    y(95) <= not(p95_out);
    p95 : perceptron
        Generic map (
            WEIGHTS => "10001",
            SHIFT => 5,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p95_in,
            y(0) => p95_out,
            y(1 to 13 - 1) => dummy95
        );


    p96_in <= x(25) & x(43) & x(77) & x(232) & x(240);
    y(96) <= not(p96_out);
    p96 : perceptron
        Generic map (
            WEIGHTS => "01110",
            SHIFT => 5,
            B => 5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p96_in,
            y(0) => p96_out,
            y(1 to 13 - 1) => dummy96
        );


    p97_in <= x(54) & x(114) & x(153) & x(229) & x(254);
    y(97) <= not(p97_out);
    p97 : perceptron
        Generic map (
            WEIGHTS => "11001",
            SHIFT => 5,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p97_in,
            y(0) => p97_out,
            y(1 to 13 - 1) => dummy97
        );


    p98_in <= x(153) & x(208) & x(223) & x(239) & x(243);
    y(98) <= not(p98_out);
    p98 : perceptron
        Generic map (
            WEIGHTS => "10101",
            SHIFT => 6,
            B => 10,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p98_in,
            y(0) => p98_out,
            y(1 to 14 - 1) => dummy98
        );


    p99_in <= x(3) & x(9) & x(34) & x(49);
    y(99) <= not(p99_out);
    p99 : perceptron
        Generic map (
            WEIGHTS => "0000",
            SHIFT => 5,
            B => -8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p99_in,
            y(0) => p99_out,
            y(1 to 12 - 1) => dummy99
        );


    p100_in <= x(30) & x(34) & x(43) & x(59) & x(84) & x(248) & x(254);
    y(100) <= not(p100_out);
    p100 : perceptron
        Generic map (
            WEIGHTS => "0100011",
            SHIFT => 5,
            B => -11,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p100_in,
            y(0) => p100_out,
            y(1 to 13 - 1) => dummy100
        );


    p101_in <= x(149) & x(254);
    y(101) <= not(p101_out);
    p101 : perceptron
        Generic map (
            WEIGHTS => "00",
            SHIFT => 6,
            B => 18,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p101_in,
            y(0) => p101_out,
            y(1 to 12 - 1) => dummy101
        );


    p102_in <= x(26) & x(41) & x(61) & x(89) & x(101) & x(104) & x(115) & x(190) & x(208) & x(229) & x(241) & x(243);
    y(102) <= not(p102_out);
    p102 : perceptron
        Generic map (
            WEIGHTS => "010001100111",
            SHIFT => 4,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p102_in,
            y(0) => p102_out,
            y(1 to 13 - 1) => dummy102
        );


    p103_in <= x(36) & x(121) & x(237);
    y(103) <= not(p103_out);
    p103 : perceptron
        Generic map (
            WEIGHTS => "011",
            SHIFT => 5,
            B => -9,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p103_in,
            y(0) => p103_out,
            y(1 to 12 - 1) => dummy103
        );


    p104_in <= x(80) & x(104) & x(153) & x(196) & x(241);
    y(104) <= not(p104_out);
    p104 : perceptron
        Generic map (
            WEIGHTS => "10100",
            SHIFT => 5,
            B => -16,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p104_in,
            y(0) => p104_out,
            y(1 to 13 - 1) => dummy104
        );


    p105_in <= x(35) & x(61) & x(78) & x(127) & x(131) & x(154) & x(155) & x(253);
    y(105) <= not(p105_out);
    p105 : perceptron
        Generic map (
            WEIGHTS => "11101100",
            SHIFT => 5,
            B => -9,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p105_in,
            y(0) => p105_out,
            y(1 to 14 - 1) => dummy105
        );


    p106_in <= x(3) & x(43) & x(77) & x(125) & x(206) & x(241);
    y(106) <= not(p106_out);
    p106 : perceptron
        Generic map (
            WEIGHTS => "111011",
            SHIFT => 5,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p106_in,
            y(0) => p106_out,
            y(1 to 13 - 1) => dummy106
        );


    p107_in <= x(66) & x(96) & x(98) & x(109) & x(125) & x(151) & x(163) & x(208);
    y(107) <= not(p107_out);
    p107 : perceptron
        Generic map (
            WEIGHTS => "11011101",
            SHIFT => 5,
            B => 5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p107_in,
            y(0) => p107_out,
            y(1 to 14 - 1) => dummy107
        );


    p108_in <= x(90) & x(101) & x(246);
    y(108) <= not(p108_out);
    p108 : perceptron
        Generic map (
            WEIGHTS => "110",
            SHIFT => 6,
            B => 10,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p108_in,
            y(0) => p108_out,
            y(1 to 13 - 1) => dummy108
        );


    p109_in <= x(43) & x(66) & x(177) & x(254);
    y(109) <= not(p109_out);
    p109 : perceptron
        Generic map (
            WEIGHTS => "0111",
            SHIFT => 6,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p109_in,
            y(0) => p109_out,
            y(1 to 13 - 1) => dummy109
        );


    p110_in <= x(109) & x(117) & x(143) & x(227) & x(248);
    y(110) <= not(p110_out);
    p110 : perceptron
        Generic map (
            WEIGHTS => "01100",
            SHIFT => 5,
            B => 17,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p110_in,
            y(0) => p110_out,
            y(1 to 13 - 1) => dummy110
        );


    p111_in <= x(65) & x(102) & x(114) & x(140) & x(216) & x(245) & x(247);
    y(111) <= not(p111_out);
    p111 : perceptron
        Generic map (
            WEIGHTS => "1110111",
            SHIFT => 5,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p111_in,
            y(0) => p111_out,
            y(1 to 13 - 1) => dummy111
        );


    p112_in(0) <= x(220);
    y(112) <= not(p112_out);
    p112 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p112_in,
            y(0) => p112_out,
            y(1 to 12 - 1) => dummy112
        );


    p113_in <= x(3) & x(7) & x(13) & x(15) & x(19) & x(35) & x(95) & x(104) & x(113) & x(240);
    y(113) <= not(p113_out);
    p113 : perceptron
        Generic map (
            WEIGHTS => "0001000100",
            SHIFT => 5,
            B => 13,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p113_in,
            y(0) => p113_out,
            y(1 to 14 - 1) => dummy113
        );


    p114_in <= x(19) & x(41) & x(69) & x(119);
    y(114) <= not(p114_out);
    p114 : perceptron
        Generic map (
            WEIGHTS => "0011",
            SHIFT => 5,
            B => 14,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p114_in,
            y(0) => p114_out,
            y(1 to 12 - 1) => dummy114
        );


    p115_in <= x(101) & x(149);
    y(115) <= not(p115_out);
    p115 : perceptron
        Generic map (
            WEIGHTS => "01",
            SHIFT => 6,
            B => -19,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p115_in,
            y(0) => p115_out,
            y(1 to 12 - 1) => dummy115
        );


    p116_in(0) <= x(241);
    y(116) <= not(p116_out);
    p116 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => -7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p116_in,
            y(0) => p116_out,
            y(1 to 12 - 1) => dummy116
        );


    p117_in <= x(15) & x(34) & x(49) & x(101) & x(104) & x(253);
    y(117) <= not(p117_out);
    p117 : perceptron
        Generic map (
            WEIGHTS => "000100",
            SHIFT => 5,
            B => 5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p117_in,
            y(0) => p117_out,
            y(1 to 13 - 1) => dummy117
        );


    p118_in <= x(66) & x(243);
    y(118) <= not(p118_out);
    p118 : perceptron
        Generic map (
            WEIGHTS => "01",
            SHIFT => 6,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p118_in,
            y(0) => p118_out,
            y(1 to 12 - 1) => dummy118
        );


    p119_in(0) <= x(143);
    y(119) <= not(p119_out);
    p119 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => 5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p119_in,
            y(0) => p119_out,
            y(1 to 12 - 1) => dummy119
        );


    p120_in <= x(3) & x(26) & x(77) & x(104) & x(121) & x(213);
    y(120) <= not(p120_out);
    p120 : perceptron
        Generic map (
            WEIGHTS => "000101",
            SHIFT => 5,
            B => 11,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p120_in,
            y(0) => p120_out,
            y(1 to 13 - 1) => dummy120
        );


    p121_in <= x(13) & x(26) & x(38) & x(115) & x(241);
    y(121) <= not(p121_out);
    p121 : perceptron
        Generic map (
            WEIGHTS => "10111",
            SHIFT => 5,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p121_in,
            y(0) => p121_out,
            y(1 to 13 - 1) => dummy121
        );


    p122_in <= x(43) & x(58) & x(66) & x(68) & x(122) & x(143) & x(157) & x(191) & x(227) & x(235) & x(248) & x(254);
    y(122) <= not(p122_out);
    p122 : perceptron
        Generic map (
            WEIGHTS => "100101010100",
            SHIFT => 4,
            B => 4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p122_in,
            y(0) => p122_out,
            y(1 to 13 - 1) => dummy122
        );


    p123_in <= x(43) & x(191) & x(235) & x(254);
    y(123) <= not(p123_out);
    p123 : perceptron
        Generic map (
            WEIGHTS => "1110",
            SHIFT => 6,
            B => 4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p123_in,
            y(0) => p123_out,
            y(1 to 14 - 1) => dummy123
        );


    p124_in <= x(81) & x(104) & x(115) & x(124) & x(229) & x(232) & x(241) & x(254);
    y(124) <= not(p124_out);
    p124 : perceptron
        Generic map (
            WEIGHTS => "11101110",
            SHIFT => 5,
            B => 4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p124_in,
            y(0) => p124_out,
            y(1 to 14 - 1) => dummy124
        );


    p125_in(0) <= x(178);
    y(125) <= not(p125_out);
    p125 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => 16,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p125_in,
            y(0) => p125_out,
            y(1 to 12 - 1) => dummy125
        );


    p126_in <= x(46) & x(51) & x(167) & x(254);
    y(126) <= not(p126_out);
    p126 : perceptron
        Generic map (
            WEIGHTS => "0001",
            SHIFT => 6,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p126_in,
            y(0) => p126_out,
            y(1 to 13 - 1) => dummy126
        );


    p127_in <= x(114) & x(129) & x(190) & x(251) & x(254);
    y(127) <= not(p127_out);
    p127 : perceptron
        Generic map (
            WEIGHTS => "10011",
            SHIFT => 5,
            B => -8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p127_in,
            y(0) => p127_out,
            y(1 to 13 - 1) => dummy127
        );


    p128_in <= x(13) & x(29) & x(49) & x(121);
    y(128) <= not(p128_out);
    p128 : perceptron
        Generic map (
            WEIGHTS => "0111",
            SHIFT => 6,
            B => -7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p128_in,
            y(0) => p128_out,
            y(1 to 13 - 1) => dummy128
        );


    p129_in <= x(101) & x(104) & x(121) & x(153) & x(155) & x(160) & x(164) & x(237);
    y(129) <= not(p129_out);
    p129 : perceptron
        Generic map (
            WEIGHTS => "01111001",
            SHIFT => 4,
            B => -7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p129_in,
            y(0) => p129_out,
            y(1 to 13 - 1) => dummy129
        );


    p130_in <= x(5) & x(48) & x(103) & x(151);
    y(130) <= not(p130_out);
    p130 : perceptron
        Generic map (
            WEIGHTS => "1111",
            SHIFT => 5,
            B => 6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p130_in,
            y(0) => p130_out,
            y(1 to 12 - 1) => dummy130
        );


    p131_in <= x(49) & x(131) & x(232);
    y(131) <= not(p131_out);
    p131 : perceptron
        Generic map (
            WEIGHTS => "010",
            SHIFT => 6,
            B => 4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p131_in,
            y(0) => p131_out,
            y(1 to 13 - 1) => dummy131
        );


    p132_in <= x(79) & x(104) & x(181);
    y(132) <= not(p132_out);
    p132 : perceptron
        Generic map (
            WEIGHTS => "101",
            SHIFT => 6,
            B => -10,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p132_in,
            y(0) => p132_out,
            y(1 to 13 - 1) => dummy132
        );


    p133_in <= x(26) & x(74) & x(76) & x(232) & x(243);
    y(133) <= not(p133_out);
    p133 : perceptron
        Generic map (
            WEIGHTS => "10000",
            SHIFT => 5,
            B => -8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p133_in,
            y(0) => p133_out,
            y(1 to 13 - 1) => dummy133
        );


    p134_in <= x(36) & x(41) & x(88) & x(91) & x(162) & x(170) & x(202);
    y(134) <= not(p134_out);
    p134 : perceptron
        Generic map (
            WEIGHTS => "0011010",
            SHIFT => 5,
            B => 4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p134_in,
            y(0) => p134_out,
            y(1 to 13 - 1) => dummy134
        );


    p135_in <= x(114) & x(232) & x(254);
    y(135) <= not(p135_out);
    p135 : perceptron
        Generic map (
            WEIGHTS => "101",
            SHIFT => 6,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p135_in,
            y(0) => p135_out,
            y(1 to 13 - 1) => dummy135
        );


    p136_in <= x(34) & x(106) & x(114) & x(179) & x(215) & x(229) & x(232) & x(241);
    y(136) <= not(p136_out);
    p136 : perceptron
        Generic map (
            WEIGHTS => "01001111",
            SHIFT => 5,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p136_in,
            y(0) => p136_out,
            y(1 to 14 - 1) => dummy136
        );


    p137_in <= x(1) & x(117) & x(124) & x(215);
    y(137) <= not(p137_out);
    p137 : perceptron
        Generic map (
            WEIGHTS => "1001",
            SHIFT => 5,
            B => -12,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p137_in,
            y(0) => p137_out,
            y(1 to 12 - 1) => dummy137
        );


    p138_in <= x(12) & x(26) & x(104) & x(115) & x(229);
    y(138) <= not(p138_out);
    p138 : perceptron
        Generic map (
            WEIGHTS => "01000",
            SHIFT => 5,
            B => -11,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p138_in,
            y(0) => p138_out,
            y(1 to 13 - 1) => dummy138
        );


    p139_in <= x(3) & x(101) & x(174) & x(215) & x(232);
    y(139) <= not(p139_out);
    p139 : perceptron
        Generic map (
            WEIGHTS => "01000",
            SHIFT => 5,
            B => 8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p139_in,
            y(0) => p139_out,
            y(1 to 13 - 1) => dummy139
        );


    p140_in <= x(86) & x(229) & x(230) & x(244);
    y(140) <= not(p140_out);
    p140 : perceptron
        Generic map (
            WEIGHTS => "0111",
            SHIFT => 5,
            B => 21,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p140_in,
            y(0) => p140_out,
            y(1 to 13 - 1) => dummy140
        );


    p141_in <= x(34) & x(43) & x(49) & x(101) & x(170) & x(210) & x(248) & x(253);
    y(141) <= not(p141_out);
    p141 : perceptron
        Generic map (
            WEIGHTS => "01010100",
            SHIFT => 5,
            B => 16,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p141_in,
            y(0) => p141_out,
            y(1 to 14 - 1) => dummy141
        );


    p142_in <= x(157) & x(241);
    y(142) <= not(p142_out);
    p142 : perceptron
        Generic map (
            WEIGHTS => "10",
            SHIFT => 6,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p142_in,
            y(0) => p142_out,
            y(1 to 12 - 1) => dummy142
        );


    p143_in <= x(26) & x(38) & x(104) & x(113) & x(115) & x(213) & x(241) & x(243);
    y(143) <= not(p143_out);
    p143 : perceptron
        Generic map (
            WEIGHTS => "01111111",
            SHIFT => 4,
            B => 7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p143_in,
            y(0) => p143_out,
            y(1 to 13 - 1) => dummy143
        );


    p144_in <= x(13) & x(33) & x(159) & x(191) & x(235) & x(248) & x(254);
    y(144) <= not(p144_out);
    p144 : perceptron
        Generic map (
            WEIGHTS => "1100011",
            SHIFT => 5,
            B => -10,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p144_in,
            y(0) => p144_out,
            y(1 to 13 - 1) => dummy144
        );


    p145_in <= x(104) & x(241);
    y(145) <= not(p145_out);
    p145 : perceptron
        Generic map (
            WEIGHTS => "00",
            SHIFT => 6,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p145_in,
            y(0) => p145_out,
            y(1 to 12 - 1) => dummy145
        );


    p146_in <= x(43) & x(230) & x(235) & x(254);
    y(146) <= not(p146_out);
    p146 : perceptron
        Generic map (
            WEIGHTS => "1110",
            SHIFT => 6,
            B => 10,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p146_in,
            y(0) => p146_out,
            y(1 to 14 - 1) => dummy146
        );


    p147_in <= x(30) & x(43) & x(59) & x(66) & x(121) & x(125) & x(164) & x(210);
    y(147) <= not(p147_out);
    p147 : perceptron
        Generic map (
            WEIGHTS => "11100110",
            SHIFT => 4,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p147_in,
            y(0) => p147_out,
            y(1 to 13 - 1) => dummy147
        );


    p148_in <= x(19) & x(41) & x(43) & x(118) & x(125) & x(170) & x(205) & x(208) & x(241);
    y(148) <= not(p148_out);
    p148 : perceptron
        Generic map (
            WEIGHTS => "111000001",
            SHIFT => 5,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p148_in,
            y(0) => p148_out,
            y(1 to 14 - 1) => dummy148
        );


    p149_in <= x(34) & x(121) & x(125) & x(153) & x(159) & x(191) & x(208) & x(248) & x(254);
    y(149) <= not(p149_out);
    p149 : perceptron
        Generic map (
            WEIGHTS => "010111000",
            SHIFT => 4,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p149_in,
            y(0) => p149_out,
            y(1 to 13 - 1) => dummy149
        );


    p150_in <= x(29) & x(106) & x(152) & x(179) & x(251);
    y(150) <= not(p150_out);
    p150 : perceptron
        Generic map (
            WEIGHTS => "00111",
            SHIFT => 5,
            B => -15,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p150_in,
            y(0) => p150_out,
            y(1 to 13 - 1) => dummy150
        );


    p151_in <= x(61) & x(114) & x(188) & x(190) & x(251) & x(254);
    y(151) <= not(p151_out);
    p151 : perceptron
        Generic map (
            WEIGHTS => "010011",
            SHIFT => 5,
            B => -7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p151_in,
            y(0) => p151_out,
            y(1 to 13 - 1) => dummy151
        );


    p152_in <= x(43) & x(77);
    y(152) <= not(p152_out);
    p152 : perceptron
        Generic map (
            WEIGHTS => "11",
            SHIFT => 6,
            B => 7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p152_in,
            y(0) => p152_out,
            y(1 to 12 - 1) => dummy152
        );


    p153_in <= x(7) & x(9) & x(49) & x(180) & x(195) & x(230);
    y(153) <= not(p153_out);
    p153 : perceptron
        Generic map (
            WEIGHTS => "100000",
            SHIFT => 5,
            B => -10,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p153_in,
            y(0) => p153_out,
            y(1 to 13 - 1) => dummy153
        );


    p154_in <= x(125) & x(153) & x(155) & x(191) & x(199) & x(208) & x(215) & x(230);
    y(154) <= not(p154_out);
    p154 : perceptron
        Generic map (
            WEIGHTS => "10000101",
            SHIFT => 4,
            B => 5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p154_in,
            y(0) => p154_out,
            y(1 to 13 - 1) => dummy154
        );


    p155_in <= x(125) & x(138) & x(153) & x(155) & x(191) & x(208) & x(248);
    y(155) <= not(p155_out);
    p155 : perceptron
        Generic map (
            WEIGHTS => "1100011",
            SHIFT => 5,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p155_in,
            y(0) => p155_out,
            y(1 to 13 - 1) => dummy155
        );


    p156_in <= x(59) & x(125) & x(153) & x(191) & x(208) & x(215) & x(254);
    y(156) <= not(p156_out);
    p156 : perceptron
        Generic map (
            WEIGHTS => "1100101",
            SHIFT => 5,
            B => 5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p156_in,
            y(0) => p156_out,
            y(1 to 13 - 1) => dummy156
        );


    p157_in <= x(3) & x(49) & x(95) & x(130) & x(220) & x(248);
    y(157) <= not(p157_out);
    p157 : perceptron
        Generic map (
            WEIGHTS => "110101",
            SHIFT => 5,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p157_in,
            y(0) => p157_out,
            y(1 to 13 - 1) => dummy157
        );


    p158_in <= x(3) & x(30) & x(43) & x(78) & x(135) & x(154) & x(157) & x(170) & x(247);
    y(158) <= not(p158_out);
    p158 : perceptron
        Generic map (
            WEIGHTS => "100101101",
            SHIFT => 5,
            B => 4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p158_in,
            y(0) => p158_out,
            y(1 to 14 - 1) => dummy158
        );


    p159_in <= x(61) & x(106) & x(114) & x(135) & x(188) & x(190) & x(233) & x(251) & x(254);
    y(159) <= not(p159_out);
    p159 : perceptron
        Generic map (
            WEIGHTS => "001000011",
            SHIFT => 5,
            B => -10,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p159_in,
            y(0) => p159_out,
            y(1 to 14 - 1) => dummy159
        );


    p160_in <= x(68) & x(142) & x(143) & x(168);
    y(160) <= not(p160_out);
    p160 : perceptron
        Generic map (
            WEIGHTS => "1011",
            SHIFT => 5,
            B => 20,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p160_in,
            y(0) => p160_out,
            y(1 to 13 - 1) => dummy160
        );


    p161_in <= x(43) & x(68) & x(159) & x(215) & x(227) & x(248);
    y(161) <= not(p161_out);
    p161 : perceptron
        Generic map (
            WEIGHTS => "111000",
            SHIFT => 5,
            B => 6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p161_in,
            y(0) => p161_out,
            y(1 to 13 - 1) => dummy161
        );


    p162_in <= x(66) & x(68);
    y(162) <= not(p162_out);
    p162 : perceptron
        Generic map (
            WEIGHTS => "01",
            SHIFT => 6,
            B => -10,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p162_in,
            y(0) => p162_out,
            y(1 to 12 - 1) => dummy162
        );


    p163_in <= x(73) & x(106) & x(191) & x(208) & x(241) & x(251);
    y(163) <= not(p163_out);
    p163 : perceptron
        Generic map (
            WEIGHTS => "001011",
            SHIFT => 6,
            B => -14,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p163_in,
            y(0) => p163_out,
            y(1 to 14 - 1) => dummy163
        );


    p164_in <= x(30) & x(131) & x(134) & x(136);
    y(164) <= not(p164_out);
    p164 : perceptron
        Generic map (
            WEIGHTS => "1011",
            SHIFT => 5,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p164_in,
            y(0) => p164_out,
            y(1 to 13 - 1) => dummy164
        );


    p165_in <= x(3) & x(49) & x(141) & x(248);
    y(165) <= not(p165_out);
    p165 : perceptron
        Generic map (
            WEIGHTS => "1101",
            SHIFT => 5,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p165_in,
            y(0) => p165_out,
            y(1 to 12 - 1) => dummy165
        );


    p166_in <= x(50) & x(130) & x(131) & x(188);
    y(166) <= not(p166_out);
    p166 : perceptron
        Generic map (
            WEIGHTS => "0100",
            SHIFT => 5,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p166_in,
            y(0) => p166_out,
            y(1 to 13 - 1) => dummy166
        );


    p167_in <= x(38) & x(90) & x(230);
    y(167) <= not(p167_out);
    p167 : perceptron
        Generic map (
            WEIGHTS => "000",
            SHIFT => 6,
            B => -7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p167_in,
            y(0) => p167_out,
            y(1 to 13 - 1) => dummy167
        );


    p168_in <= x(30) & x(43) & x(59) & x(194) & x(254);
    y(168) <= not(p168_out);
    p168 : perceptron
        Generic map (
            WEIGHTS => "11110",
            SHIFT => 5,
            B => 13,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p168_in,
            y(0) => p168_out,
            y(1 to 13 - 1) => dummy168
        );


    p169_in <= x(43) & x(159) & x(191) & x(229) & x(230) & x(254);
    y(169) <= not(p169_out);
    p169 : perceptron
        Generic map (
            WEIGHTS => "000001",
            SHIFT => 5,
            B => -6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p169_in,
            y(0) => p169_out,
            y(1 to 13 - 1) => dummy169
        );


    p170_in <= x(49) & x(241) & x(254);
    y(170) <= not(p170_out);
    p170 : perceptron
        Generic map (
            WEIGHTS => "100",
            SHIFT => 6,
            B => -7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p170_in,
            y(0) => p170_out,
            y(1 to 13 - 1) => dummy170
        );


    p171_in <= x(36) & x(43) & x(111) & x(134);
    y(171) <= not(p171_out);
    p171 : perceptron
        Generic map (
            WEIGHTS => "0010",
            SHIFT => 6,
            B => 18,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p171_in,
            y(0) => p171_out,
            y(1 to 13 - 1) => dummy171
        );


    p172_in <= x(83) & x(114) & x(129) & x(188) & x(251);
    y(172) <= not(p172_out);
    p172 : perceptron
        Generic map (
            WEIGHTS => "10110",
            SHIFT => 5,
            B => 13,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p172_in,
            y(0) => p172_out,
            y(1 to 13 - 1) => dummy172
        );


    p173_in <= x(26) & x(43) & x(59) & x(61) & x(63);
    y(173) <= not(p173_out);
    p173 : perceptron
        Generic map (
            WEIGHTS => "10001",
            SHIFT => 5,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p173_in,
            y(0) => p173_out,
            y(1 to 13 - 1) => dummy173
        );


    p174_in <= x(32) & x(101) & x(104) & x(248) & x(253);
    y(174) <= not(p174_out);
    p174 : perceptron
        Generic map (
            WEIGHTS => "00111",
            SHIFT => 5,
            B => -11,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p174_in,
            y(0) => p174_out,
            y(1 to 13 - 1) => dummy174
        );


    p175_in <= x(36) & x(101) & x(121);
    y(175) <= not(p175_out);
    p175 : perceptron
        Generic map (
            WEIGHTS => "001",
            SHIFT => 5,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p175_in,
            y(0) => p175_out,
            y(1 to 12 - 1) => dummy175
        );


    p176_in <= x(3) & x(77) & x(157);
    y(176) <= not(p176_out);
    p176 : perceptron
        Generic map (
            WEIGHTS => "001",
            SHIFT => 6,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p176_in,
            y(0) => p176_out,
            y(1 to 13 - 1) => dummy176
        );


    p177_in <= x(106) & x(114) & x(190) & x(233) & x(251);
    y(177) <= not(p177_out);
    p177 : perceptron
        Generic map (
            WEIGHTS => "10110",
            SHIFT => 5,
            B => 8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p177_in,
            y(0) => p177_out,
            y(1 to 13 - 1) => dummy177
        );


    p178_in <= x(7) & x(43) & x(125) & x(191) & x(208) & x(230) & x(241);
    y(178) <= not(p178_out);
    p178 : perceptron
        Generic map (
            WEIGHTS => "0101011",
            SHIFT => 5,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p178_in,
            y(0) => p178_out,
            y(1 to 13 - 1) => dummy178
        );


    p179_in <= x(23) & x(57) & x(101) & x(127);
    y(179) <= not(p179_out);
    p179 : perceptron
        Generic map (
            WEIGHTS => "1110",
            SHIFT => 6,
            B => -18,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p179_in,
            y(0) => p179_out,
            y(1 to 13 - 1) => dummy179
        );


    p180_in <= x(3) & x(66) & x(77) & x(84) & x(89) & x(104) & x(153) & x(177) & x(229) & x(254);
    y(180) <= not(p180_out);
    p180 : perceptron
        Generic map (
            WEIGHTS => "1111100101",
            SHIFT => 5,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p180_in,
            y(0) => p180_out,
            y(1 to 14 - 1) => dummy180
        );


    p181_in <= x(61) & x(106) & x(114) & x(190) & x(233) & x(254);
    y(181) <= not(p181_out);
    p181 : perceptron
        Generic map (
            WEIGHTS => "110110",
            SHIFT => 5,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p181_in,
            y(0) => p181_out,
            y(1 to 13 - 1) => dummy181
        );


    p182_in <= x(15) & x(24);
    y(182) <= not(p182_out);
    p182 : perceptron
        Generic map (
            WEIGHTS => "11",
            SHIFT => 6,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p182_in,
            y(0) => p182_out,
            y(1 to 12 - 1) => dummy182
        );


    p183_in <= x(178) & x(191) & x(206);
    y(183) <= not(p183_out);
    p183 : perceptron
        Generic map (
            WEIGHTS => "000",
            SHIFT => 6,
            B => 18,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p183_in,
            y(0) => p183_out,
            y(1 to 13 - 1) => dummy183
        );


    p184_in <= x(43) & x(55) & x(80) & x(121) & x(174) & x(232);
    y(184) <= not(p184_out);
    p184 : perceptron
        Generic map (
            WEIGHTS => "111111",
            SHIFT => 5,
            B => -7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p184_in,
            y(0) => p184_out,
            y(1 to 13 - 1) => dummy184
        );


    p185_in <= x(56) & x(79) & x(152) & x(188) & x(190);
    y(185) <= not(p185_out);
    p185 : perceptron
        Generic map (
            WEIGHTS => "00100",
            SHIFT => 5,
            B => -9,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p185_in,
            y(0) => p185_out,
            y(1 to 13 - 1) => dummy185
        );


    p186_in <= x(43) & x(77) & x(90) & x(241);
    y(186) <= not(p186_out);
    p186 : perceptron
        Generic map (
            WEIGHTS => "0010",
            SHIFT => 5,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p186_in,
            y(0) => p186_out,
            y(1 to 12 - 1) => dummy186
        );


    p187_in <= x(63) & x(90) & x(101) & x(155);
    y(187) <= not(p187_out);
    p187 : perceptron
        Generic map (
            WEIGHTS => "1000",
            SHIFT => 5,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p187_in,
            y(0) => p187_out,
            y(1 to 12 - 1) => dummy187
        );


    p188_in <= x(174) & x(248);
    y(188) <= not(p188_out);
    p188 : perceptron
        Generic map (
            WEIGHTS => "00",
            SHIFT => 6,
            B => 28,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p188_in,
            y(0) => p188_out,
            y(1 to 12 - 1) => dummy188
        );


    p189_in <= x(12) & x(13) & x(26) & x(38) & x(104) & x(115) & x(190) & x(229) & x(241) & x(243);
    y(189) <= not(p189_out);
    p189 : perceptron
        Generic map (
            WEIGHTS => "1101110111",
            SHIFT => 4,
            B => 5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p189_in,
            y(0) => p189_out,
            y(1 to 13 - 1) => dummy189
        );


    p190_in <= x(74) & x(76) & x(81) & x(167) & x(232);
    y(190) <= not(p190_out);
    p190 : perceptron
        Generic map (
            WEIGHTS => "00000",
            SHIFT => 5,
            B => -11,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p190_in,
            y(0) => p190_out,
            y(1 to 13 - 1) => dummy190
        );


    p191_in <= x(13) & x(41) & x(63) & x(100) & x(115) & x(241);
    y(191) <= not(p191_out);
    p191 : perceptron
        Generic map (
            WEIGHTS => "110111",
            SHIFT => 5,
            B => -12,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p191_in,
            y(0) => p191_out,
            y(1 to 13 - 1) => dummy191
        );


    p192_in <= x(101) & x(123) & x(138) & x(230);
    y(192) <= not(p192_out);
    p192 : perceptron
        Generic map (
            WEIGHTS => "0110",
            SHIFT => 5,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p192_in,
            y(0) => p192_out,
            y(1 to 13 - 1) => dummy192
        );


    p193_in <= x(230) & x(241);
    y(193) <= not(p193_out);
    p193 : perceptron
        Generic map (
            WEIGHTS => "01",
            SHIFT => 6,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p193_in,
            y(0) => p193_out,
            y(1 to 12 - 1) => dummy193
        );


    p194_in <= x(125) & x(153) & x(191) & x(208);
    y(194) <= not(p194_out);
    p194 : perceptron
        Generic map (
            WEIGHTS => "0110",
            SHIFT => 5,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p194_in,
            y(0) => p194_out,
            y(1 to 13 - 1) => dummy194
        );


    p195_in(0) <= x(252);
    y(195) <= not(p195_out);
    p195 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p195_in,
            y(0) => p195_out,
            y(1 to 12 - 1) => dummy195
        );


    p196_in <= x(41) & x(101) & x(104) & x(115) & x(190) & x(229) & x(241) & x(253);
    y(196) <= not(p196_out);
    p196 : perceptron
        Generic map (
            WEIGHTS => "01001000",
            SHIFT => 5,
            B => 4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p196_in,
            y(0) => p196_out,
            y(1 to 14 - 1) => dummy196
        );


    p197_in <= x(7) & x(49) & x(153) & x(157);
    y(197) <= not(p197_out);
    p197 : perceptron
        Generic map (
            WEIGHTS => "1011",
            SHIFT => 5,
            B => 4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p197_in,
            y(0) => p197_out,
            y(1 to 12 - 1) => dummy197
        );


    p198_in <= x(9) & x(49) & x(232);
    y(198) <= not(p198_out);
    p198 : perceptron
        Generic map (
            WEIGHTS => "000",
            SHIFT => 6,
            B => -7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p198_in,
            y(0) => p198_out,
            y(1 to 13 - 1) => dummy198
        );


    p199_in <= x(101) & x(104) & x(121) & x(253);
    y(199) <= not(p199_out);
    p199 : perceptron
        Generic map (
            WEIGHTS => "1000",
            SHIFT => 5,
            B => 8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p199_in,
            y(0) => p199_out,
            y(1 to 13 - 1) => dummy199
        );


    p200_in <= x(34) & x(254);
    y(200) <= not(p200_out);
    p200 : perceptron
        Generic map (
            WEIGHTS => "11",
            SHIFT => 6,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p200_in,
            y(0) => p200_out,
            y(1 to 12 - 1) => dummy200
        );


    p201_in <= x(77) & x(229) & x(246);
    y(201) <= not(p201_out);
    p201 : perceptron
        Generic map (
            WEIGHTS => "100",
            SHIFT => 6,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p201_in,
            y(0) => p201_out,
            y(1 to 13 - 1) => dummy201
        );


    p202_in <= x(8) & x(96) & x(208) & x(210);
    y(202) <= not(p202_out);
    p202 : perceptron
        Generic map (
            WEIGHTS => "1001",
            SHIFT => 5,
            B => 6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p202_in,
            y(0) => p202_out,
            y(1 to 12 - 1) => dummy202
        );


    p203_in <= x(92) & x(106) & x(150);
    y(203) <= not(p203_out);
    p203 : perceptron
        Generic map (
            WEIGHTS => "100",
            SHIFT => 6,
            B => 14,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p203_in,
            y(0) => p203_out,
            y(1 to 13 - 1) => dummy203
        );


    p204_in <= x(47) & x(93) & x(101) & x(118) & x(131) & x(174) & x(230);
    y(204) <= not(p204_out);
    p204 : perceptron
        Generic map (
            WEIGHTS => "1011001",
            SHIFT => 5,
            B => 7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p204_in,
            y(0) => p204_out,
            y(1 to 13 - 1) => dummy204
        );


    p205_in <= x(43) & x(153) & x(157) & x(249);
    y(205) <= not(p205_out);
    p205 : perceptron
        Generic map (
            WEIGHTS => "1001",
            SHIFT => 5,
            B => 4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p205_in,
            y(0) => p205_out,
            y(1 to 13 - 1) => dummy205
        );


    p206_in <= x(13) & x(58) & x(68) & x(141) & x(159) & x(191) & x(227) & x(248);
    y(206) <= not(p206_out);
    p206 : perceptron
        Generic map (
            WEIGHTS => "00111100",
            SHIFT => 4,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p206_in,
            y(0) => p206_out,
            y(1 to 13 - 1) => dummy206
        );


    p207_in <= x(3) & x(77) & x(86) & x(121) & x(125) & x(177) & x(208);
    y(207) <= not(p207_out);
    p207 : perceptron
        Generic map (
            WEIGHTS => "0010101",
            SHIFT => 5,
            B => -10,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p207_in,
            y(0) => p207_out,
            y(1 to 13 - 1) => dummy207
        );


    p208_in <= x(3) & x(41);
    y(208) <= not(p208_out);
    p208 : perceptron
        Generic map (
            WEIGHTS => "11",
            SHIFT => 6,
            B => -17,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p208_in,
            y(0) => p208_out,
            y(1 to 12 - 1) => dummy208
        );


    p209_in <= x(7) & x(13) & x(43) & x(58) & x(66) & x(68) & x(86) & x(141) & x(159) & x(178) & x(191);
    y(209) <= not(p209_out);
    p209 : perceptron
        Generic map (
            WEIGHTS => "00100101111",
            SHIFT => 4,
            B => -7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p209_in,
            y(0) => p209_out,
            y(1 to 13 - 1) => dummy209
        );


    p210_in <= x(13) & x(59) & x(153) & x(191);
    y(210) <= not(p210_out);
    p210 : perceptron
        Generic map (
            WEIGHTS => "1100",
            SHIFT => 5,
            B => 11,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p210_in,
            y(0) => p210_out,
            y(1 to 12 - 1) => dummy210
        );


    p211_in <= x(153) & x(208) & x(229);
    y(211) <= not(p211_out);
    p211 : perceptron
        Generic map (
            WEIGHTS => "010",
            SHIFT => 6,
            B => -9,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p211_in,
            y(0) => p211_out,
            y(1 to 13 - 1) => dummy211
        );


    p212_in <= x(168) & x(170) & x(237);
    y(212) <= not(p212_out);
    p212 : perceptron
        Generic map (
            WEIGHTS => "011",
            SHIFT => 6,
            B => -45,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p212_in,
            y(0) => p212_out,
            y(1 to 13 - 1) => dummy212
        );


    p213_in <= x(22) & x(68) & x(190);
    y(213) <= not(p213_out);
    p213 : perceptron
        Generic map (
            WEIGHTS => "000",
            SHIFT => 6,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p213_in,
            y(0) => p213_out,
            y(1 to 13 - 1) => dummy213
        );


    p214_in <= x(14) & x(25) & x(124) & x(208);
    y(214) <= not(p214_out);
    p214 : perceptron
        Generic map (
            WEIGHTS => "0011",
            SHIFT => 6,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p214_in,
            y(0) => p214_out,
            y(1 to 13 - 1) => dummy214
        );


    p215_in <= x(34) & x(79) & x(89) & x(153) & x(191) & x(229);
    y(215) <= not(p215_out);
    p215 : perceptron
        Generic map (
            WEIGHTS => "000111",
            SHIFT => 5,
            B => -6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p215_in,
            y(0) => p215_out,
            y(1 to 13 - 1) => dummy215
        );


    p216_in <= x(80) & x(121) & x(123) & x(178);
    y(216) <= not(p216_out);
    p216 : perceptron
        Generic map (
            WEIGHTS => "0010",
            SHIFT => 6,
            B => 10,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p216_in,
            y(0) => p216_out,
            y(1 to 14 - 1) => dummy216
        );


    p217_in <= x(1) & x(90) & x(117) & x(220);
    y(217) <= not(p217_out);
    p217 : perceptron
        Generic map (
            WEIGHTS => "1101",
            SHIFT => 5,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p217_in,
            y(0) => p217_out,
            y(1 to 12 - 1) => dummy217
        );


    p218_in <= x(3) & x(7) & x(24) & x(49) & x(206) & x(246);
    y(218) <= not(p218_out);
    p218 : perceptron
        Generic map (
            WEIGHTS => "010000",
            SHIFT => 5,
            B => 4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p218_in,
            y(0) => p218_out,
            y(1 to 13 - 1) => dummy218
        );


    p219_in <= x(43) & x(115) & x(149) & x(241) & x(243);
    y(219) <= not(p219_out);
    p219 : perceptron
        Generic map (
            WEIGHTS => "11011",
            SHIFT => 5,
            B => 9,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p219_in,
            y(0) => p219_out,
            y(1 to 13 - 1) => dummy219
        );


    p220_in <= x(59) & x(68) & x(121) & x(124) & x(125) & x(153) & x(155) & x(199) & x(215) & x(230);
    y(220) <= not(p220_out);
    p220 : perceptron
        Generic map (
            WEIGHTS => "0010011110",
            SHIFT => 4,
            B => -9,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p220_in,
            y(0) => p220_out,
            y(1 to 13 - 1) => dummy220
        );


    p222_in <= x(1) & x(114) & x(131);
    y(222) <= not(p222_out);
    p222 : perceptron
        Generic map (
            WEIGHTS => "101",
            SHIFT => 6,
            B => 5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p222_in,
            y(0) => p222_out,
            y(1 to 13 - 1) => dummy222
        );


    p223_in <= x(43) & x(59) & x(104) & x(121) & x(164);
    y(223) <= not(p223_out);
    p223 : perceptron
        Generic map (
            WEIGHTS => "11001",
            SHIFT => 5,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p223_in,
            y(0) => p223_out,
            y(1 to 13 - 1) => dummy223
        );


    p224_in <= x(13) & x(66) & x(68) & x(141) & x(143) & x(157) & x(159) & x(227) & x(248);
    y(224) <= not(p224_out);
    p224 : perceptron
        Generic map (
            WEIGHTS => "001110100",
            SHIFT => 4,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p224_in,
            y(0) => p224_out,
            y(1 to 13 - 1) => dummy224
        );


    p225_in <= x(3) & x(157) & x(248);
    y(225) <= not(p225_out);
    p225 : perceptron
        Generic map (
            WEIGHTS => "011",
            SHIFT => 6,
            B => -11,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p225_in,
            y(0) => p225_out,
            y(1 to 13 - 1) => dummy225
        );


    p226_in <= x(10) & x(29) & x(31) & x(114) & x(120) & x(135) & x(137) & x(152) & x(190) & x(251);
    y(226) <= not(p226_out);
    p226 : perceptron
        Generic map (
            WEIGHTS => "0011000101",
            SHIFT => 4,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p226_in,
            y(0) => p226_out,
            y(1 to 13 - 1) => dummy226
        );


    p227_in <= x(77) & x(121) & x(157);
    y(227) <= not(p227_out);
    p227 : perceptron
        Generic map (
            WEIGHTS => "110",
            SHIFT => 6,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p227_in,
            y(0) => p227_out,
            y(1 to 13 - 1) => dummy227
        );


    p228_in <= x(34) & x(59) & x(101) & x(141) & x(208) & x(227) & x(248);
    y(228) <= not(p228_out);
    p228 : perceptron
        Generic map (
            WEIGHTS => "0111000",
            SHIFT => 5,
            B => 9,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p228_in,
            y(0) => p228_out,
            y(1 to 13 - 1) => dummy228
        );


    p229_in <= x(49) & x(90) & x(153) & x(203) & x(220);
    y(229) <= not(p229_out);
    p229 : perceptron
        Generic map (
            WEIGHTS => "10010",
            SHIFT => 5,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p229_in,
            y(0) => p229_out,
            y(1 to 13 - 1) => dummy229
        );


    p230_in <= x(93) & x(157) & x(250);
    y(230) <= not(p230_out);
    p230 : perceptron
        Generic map (
            WEIGHTS => "011",
            SHIFT => 6,
            B => 30,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p230_in,
            y(0) => p230_out,
            y(1 to 13 - 1) => dummy230
        );


    p231_in <= x(78) & x(121) & x(143) & x(227) & x(248);
    y(231) <= not(p231_out);
    p231 : perceptron
        Generic map (
            WEIGHTS => "01100",
            SHIFT => 5,
            B => 11,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p231_in,
            y(0) => p231_out,
            y(1 to 13 - 1) => dummy231
        );


    p232_in <= x(41) & x(75) & x(118) & x(154) & x(190) & x(192) & x(237) & x(241);
    y(232) <= not(p232_out);
    p232 : perceptron
        Generic map (
            WEIGHTS => "11110011",
            SHIFT => 5,
            B => -15,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p232_in,
            y(0) => p232_out,
            y(1 to 14 - 1) => dummy232
        );


    p233_in <= x(43) & x(191) & x(254);
    y(233) <= not(p233_out);
    p233 : perceptron
        Generic map (
            WEIGHTS => "110",
            SHIFT => 6,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p233_in,
            y(0) => p233_out,
            y(1 to 13 - 1) => dummy233
        );


    p234_in <= x(66) & x(143);
    y(234) <= not(p234_out);
    p234 : perceptron
        Generic map (
            WEIGHTS => "01",
            SHIFT => 6,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p234_in,
            y(0) => p234_out,
            y(1 to 12 - 1) => dummy234
        );


    p235_in <= x(7) & x(49) & x(81) & x(131) & x(135) & x(187) & x(230) & x(232);
    y(235) <= not(p235_out);
    p235 : perceptron
        Generic map (
            WEIGHTS => "10010100",
            SHIFT => 5,
            B => 4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p235_in,
            y(0) => p235_out,
            y(1 to 14 - 1) => dummy235
        );


    p236_in <= x(39) & x(77) & x(79) & x(81) & x(89) & x(92) & x(129) & x(177) & x(205);
    y(236) <= not(p236_out);
    p236 : perceptron
        Generic map (
            WEIGHTS => "100101101",
            SHIFT => 5,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p236_in,
            y(0) => p236_out,
            y(1 to 14 - 1) => dummy236
        );


    p237_in <= x(191) & x(214);
    y(237) <= not(p237_out);
    p237 : perceptron
        Generic map (
            WEIGHTS => "10",
            SHIFT => 6,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p237_in,
            y(0) => p237_out,
            y(1 to 12 - 1) => dummy237
        );


    p238_in <= x(25) & x(34) & x(110) & x(114) & x(128) & x(191) & x(203) & x(208) & x(254);
    y(238) <= not(p238_out);
    p238 : perceptron
        Generic map (
            WEIGHTS => "010100011",
            SHIFT => 5,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p238_in,
            y(0) => p238_out,
            y(1 to 14 - 1) => dummy238
        );


    p239_in <= x(66) & x(86) & x(89) & x(194) & x(246) & x(254);
    y(239) <= not(p239_out);
    p239 : perceptron
        Generic map (
            WEIGHTS => "010110",
            SHIFT => 5,
            B => 4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p239_in,
            y(0) => p239_out,
            y(1 to 13 - 1) => dummy239
        );


    p240_in <= x(3) & x(66) & x(248);
    y(240) <= not(p240_out);
    p240 : perceptron
        Generic map (
            WEIGHTS => "000",
            SHIFT => 5,
            B => 10,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p240_in,
            y(0) => p240_out,
            y(1 to 12 - 1) => dummy240
        );


    p241_in <= x(131) & x(232);
    y(241) <= not(p241_out);
    p241 : perceptron
        Generic map (
            WEIGHTS => "01",
            SHIFT => 6,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p241_in,
            y(0) => p241_out,
            y(1 to 12 - 1) => dummy241
        );


    p242_in <= x(79) & x(114) & x(135) & x(150) & x(152) & x(159) & x(181) & x(190) & x(251);
    y(242) <= not(p242_out);
    p242 : perceptron
        Generic map (
            WEIGHTS => "010010001",
            SHIFT => 5,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p242_in,
            y(0) => p242_out,
            y(1 to 14 - 1) => dummy242
        );


    p243_in <= x(15) & x(25) & x(37) & x(129) & x(222);
    y(243) <= not(p243_out);
    p243 : perceptron
        Generic map (
            WEIGHTS => "01010",
            SHIFT => 5,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p243_in,
            y(0) => p243_out,
            y(1 to 13 - 1) => dummy243
        );


    p244_in <= x(15) & x(153) & x(208) & x(223) & x(239) & x(243);
    y(244) <= not(p244_out);
    p244 : perceptron
        Generic map (
            WEIGHTS => "101010",
            SHIFT => 5,
            B => -8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p244_in,
            y(0) => p244_out,
            y(1 to 13 - 1) => dummy244
        );


    p246_in <= x(61) & x(114);
    y(246) <= not(p246_out);
    p246 : perceptron
        Generic map (
            WEIGHTS => "10",
            SHIFT => 6,
            B => -13,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p246_in,
            y(0) => p246_out,
            y(1 to 12 - 1) => dummy246
        );


    p247_in(0) <= x(66);
    y(247) <= not(p247_out);
    p247 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p247_in,
            y(0) => p247_out,
            y(1 to 12 - 1) => dummy247
        );


    p248_in <= x(3) & x(5) & x(32) & x(34) & x(43) & x(77) & x(104) & x(248) & x(253);
    y(248) <= not(p248_out);
    p248 : perceptron
        Generic map (
            WEIGHTS => "101011000",
            SHIFT => 5,
            B => 7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p248_in,
            y(0) => p248_out,
            y(1 to 14 - 1) => dummy248
        );


    p249_in <= x(15) & x(46) & x(109) & x(157) & x(162) & x(203);
    y(249) <= not(p249_out);
    p249 : perceptron
        Generic map (
            WEIGHTS => "011110",
            SHIFT => 5,
            B => -7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p249_in,
            y(0) => p249_out,
            y(1 to 13 - 1) => dummy249
        );


    p250_in <= x(4) & x(5) & x(36) & x(43) & x(63) & x(80) & x(93) & x(129) & x(134) & x(157) & x(159) & x(235) & x(254) & x(255);
    y(250) <= not(p250_out);
    p250 : perceptron
        Generic map (
            WEIGHTS => "11000001010011",
            SHIFT => 4,
            B => 6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p250_in,
            y(0) => p250_out,
            y(1 to 13 - 1) => dummy250
        );


    p251_in <= x(3) & x(43) & x(177) & x(205);
    y(251) <= not(p251_out);
    p251 : perceptron
        Generic map (
            WEIGHTS => "1110",
            SHIFT => 5,
            B => 5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p251_in,
            y(0) => p251_out,
            y(1 to 12 - 1) => dummy251
        );


    p252_in <= x(58) & x(131) & x(194) & x(235) & x(254);
    y(252) <= not(p252_out);
    p252 : perceptron
        Generic map (
            WEIGHTS => "11001",
            SHIFT => 5,
            B => -17,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p252_in,
            y(0) => p252_out,
            y(1 to 13 - 1) => dummy252
        );


    p253_in <= x(22) & x(106) & x(114) & x(135) & x(179) & x(190) & x(251) & x(254);
    y(253) <= not(p253_out);
    p253 : perceptron
        Generic map (
            WEIGHTS => "11010100",
            SHIFT => 5,
            B => 8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p253_in,
            y(0) => p253_out,
            y(1 to 14 - 1) => dummy253
        );


    p254_in <= x(43) & x(68) & x(101) & x(104) & x(121) & x(124) & x(164) & x(230) & x(237);
    y(254) <= not(p254_out);
    p254 : perceptron
        Generic map (
            WEIGHTS => "000110001",
            SHIFT => 5,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p254_in,
            y(0) => p254_out,
            y(1 to 14 - 1) => dummy254
        );


    p255_in <= x(6) & x(8) & x(15) & x(86) & x(230);
    y(255) <= not(p255_out);
    p255 : perceptron
        Generic map (
            WEIGHTS => "11101",
            SHIFT => 5,
            B => 4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p255_in,
            y(0) => p255_out,
            y(1 to 13 - 1) => dummy255
        );



end layer_3;

architecture layer_4 of layer is

    Component perceptron
    Generic (
        WEIGHTS : STD_LOGIC_VECTOR := (others => '0');
        SHIFT : Integer;     -- number of shift (left + or right -)
        B : Integer;          -- bias of batch norm
        BATCH_POSITIVE : Boolean    
    );
    Port ( 
        x : in STD_LOGIC_VECTOR;
        y : out STD_LOGIC_VECTOR
   );
    end component;
    
    -- Signals
    signal p0_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p0_out : STD_LOGIC;
	signal p1_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p1_out : STD_LOGIC;
	signal p2_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p2_out : STD_LOGIC;
	signal p3_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p3_out : STD_LOGIC;
	signal p4_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p4_out : STD_LOGIC;
	signal p5_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p5_out : STD_LOGIC;
	signal p6_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p6_out : STD_LOGIC;
	signal p7_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p7_out : STD_LOGIC;
	signal p8_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p8_out : STD_LOGIC;
	signal p9_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p9_out : STD_LOGIC;
	signal p10_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p10_out : STD_LOGIC;
	signal p11_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p11_out : STD_LOGIC;
	signal p12_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p12_out : STD_LOGIC;
	signal p13_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p13_out : STD_LOGIC;
	signal p14_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p14_out : STD_LOGIC;
	signal p15_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p15_out : STD_LOGIC;
	signal p16_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p16_out : STD_LOGIC;
	signal p17_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p17_out : STD_LOGIC;
	signal p18_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p18_out : STD_LOGIC;
	signal p19_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p19_out : STD_LOGIC;
	signal p20_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p20_out : STD_LOGIC;
	signal p21_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p21_out : STD_LOGIC;
	signal p22_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p22_out : STD_LOGIC;
	signal p23_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p23_out : STD_LOGIC;
	signal p24_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p24_out : STD_LOGIC;
	signal p25_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p25_out : STD_LOGIC;
	signal p26_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p26_out : STD_LOGIC;
	signal p27_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p27_out : STD_LOGIC;
	signal p28_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p28_out : STD_LOGIC;
	signal p29_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p29_out : STD_LOGIC;
	signal p30_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p30_out : STD_LOGIC;
	signal p31_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p31_out : STD_LOGIC;
	signal p32_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p32_out : STD_LOGIC;
	signal p33_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p33_out : STD_LOGIC;
	signal p34_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p34_out : STD_LOGIC;
	signal p35_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p35_out : STD_LOGIC;
	signal p36_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p36_out : STD_LOGIC;
	signal p37_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p37_out : STD_LOGIC;
	signal p38_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p38_out : STD_LOGIC;
	signal p39_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p39_out : STD_LOGIC;
	signal p40_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p40_out : STD_LOGIC;
	signal p41_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p41_out : STD_LOGIC;
	signal p42_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p42_out : STD_LOGIC;
	signal p43_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p43_out : STD_LOGIC;
	signal p44_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p44_out : STD_LOGIC;
	signal p45_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p45_out : STD_LOGIC;
	signal p46_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p46_out : STD_LOGIC;
	signal p47_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p47_out : STD_LOGIC;
	signal p48_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p48_out : STD_LOGIC;
	signal p49_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p49_out : STD_LOGIC;
	signal p50_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p50_out : STD_LOGIC;
	signal p51_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p51_out : STD_LOGIC;
	signal p52_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p52_out : STD_LOGIC;
	signal p53_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p53_out : STD_LOGIC;
	signal p54_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p54_out : STD_LOGIC;
	signal p55_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p55_out : STD_LOGIC;
	signal p56_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p56_out : STD_LOGIC;
	signal p57_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p57_out : STD_LOGIC;
	signal p58_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p58_out : STD_LOGIC;
	signal p59_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p59_out : STD_LOGIC;
	signal p60_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p60_out : STD_LOGIC;
	signal p61_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p61_out : STD_LOGIC;
	signal p62_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p62_out : STD_LOGIC;
	signal p63_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p63_out : STD_LOGIC;
	signal p64_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p64_out : STD_LOGIC;
	signal p65_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p65_out : STD_LOGIC;
	signal p66_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p66_out : STD_LOGIC;
	signal p67_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p67_out : STD_LOGIC;
	signal p68_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p68_out : STD_LOGIC;
	signal p69_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p69_out : STD_LOGIC;
	signal p70_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p70_out : STD_LOGIC;
	signal p71_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p71_out : STD_LOGIC;
	signal p72_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p72_out : STD_LOGIC;
	signal p73_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p73_out : STD_LOGIC;
	signal p74_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p74_out : STD_LOGIC;
	signal p75_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p75_out : STD_LOGIC;
	signal p76_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p76_out : STD_LOGIC;
	signal p77_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p77_out : STD_LOGIC;
	signal p78_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p78_out : STD_LOGIC;
	signal p79_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p79_out : STD_LOGIC;
	signal p80_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p80_out : STD_LOGIC;
	signal p81_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p81_out : STD_LOGIC;
	signal p82_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p82_out : STD_LOGIC;
	signal p83_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p83_out : STD_LOGIC;
	signal p84_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p84_out : STD_LOGIC;
	signal p85_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p85_out : STD_LOGIC;
	signal p86_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p86_out : STD_LOGIC;
	signal p87_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p87_out : STD_LOGIC;
	signal p88_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p88_out : STD_LOGIC;
	signal p89_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p89_out : STD_LOGIC;
	signal p90_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p90_out : STD_LOGIC;
	signal p91_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p91_out : STD_LOGIC;
	signal p92_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p92_out : STD_LOGIC;
	signal p93_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p93_out : STD_LOGIC;
	signal p94_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p94_out : STD_LOGIC;
	signal p95_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p95_out : STD_LOGIC;
	signal p96_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p96_out : STD_LOGIC;
	signal p97_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p97_out : STD_LOGIC;
	signal p98_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p98_out : STD_LOGIC;
	signal p99_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p99_out : STD_LOGIC;
	signal p100_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p100_out : STD_LOGIC;
	signal p101_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p101_out : STD_LOGIC;
	signal p102_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p102_out : STD_LOGIC;
	signal p103_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p103_out : STD_LOGIC;
	signal p104_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p104_out : STD_LOGIC;
	signal p105_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p105_out : STD_LOGIC;
	signal p106_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p106_out : STD_LOGIC;
	signal p107_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p107_out : STD_LOGIC;
	signal p108_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p108_out : STD_LOGIC;
	signal p109_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p109_out : STD_LOGIC;
	signal p110_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p110_out : STD_LOGIC;
	signal p111_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p111_out : STD_LOGIC;
	signal p112_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p112_out : STD_LOGIC;
	signal p113_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p113_out : STD_LOGIC;
	signal p114_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p114_out : STD_LOGIC;
	signal p115_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p115_out : STD_LOGIC;
	signal p116_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p116_out : STD_LOGIC;
	signal p117_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p117_out : STD_LOGIC;
	signal p118_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p118_out : STD_LOGIC;
	signal p119_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p119_out : STD_LOGIC;
	signal p120_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p120_out : STD_LOGIC;
	signal p121_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p121_out : STD_LOGIC;
	signal p122_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p122_out : STD_LOGIC;
	signal p123_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p123_out : STD_LOGIC;
	signal p124_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p124_out : STD_LOGIC;
	signal p125_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p125_out : STD_LOGIC;
	signal p126_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p126_out : STD_LOGIC;
	signal p127_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p127_out : STD_LOGIC;
	signal p128_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p128_out : STD_LOGIC;
	signal p129_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p129_out : STD_LOGIC;
	signal p130_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p130_out : STD_LOGIC;
	signal p131_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p131_out : STD_LOGIC;
	signal p132_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p132_out : STD_LOGIC;
	signal p133_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p133_out : STD_LOGIC;
	signal p134_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p134_out : STD_LOGIC;
	signal p135_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p135_out : STD_LOGIC;
	signal p136_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p136_out : STD_LOGIC;
	signal p137_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p137_out : STD_LOGIC;
	signal p138_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p138_out : STD_LOGIC;
	signal p139_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p139_out : STD_LOGIC;
	signal p140_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p140_out : STD_LOGIC;
	signal p141_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p141_out : STD_LOGIC;
	signal p142_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p142_out : STD_LOGIC;
	signal p143_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p143_out : STD_LOGIC;
	signal p144_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p144_out : STD_LOGIC;
	signal p145_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p145_out : STD_LOGIC;
	signal p146_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p146_out : STD_LOGIC;
	signal p147_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p147_out : STD_LOGIC;
	signal p148_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p148_out : STD_LOGIC;
	signal p149_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p149_out : STD_LOGIC;
	signal p150_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p150_out : STD_LOGIC;
	signal p151_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p151_out : STD_LOGIC;
	signal p152_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p152_out : STD_LOGIC;
	signal p153_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p153_out : STD_LOGIC;
	signal p154_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p154_out : STD_LOGIC;
	signal p155_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p155_out : STD_LOGIC;
	signal p156_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p156_out : STD_LOGIC;
	signal p157_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p157_out : STD_LOGIC;
	signal p158_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p158_out : STD_LOGIC;
	signal p159_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p159_out : STD_LOGIC;
	signal p160_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p160_out : STD_LOGIC;
	signal p161_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p161_out : STD_LOGIC;
	signal p162_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p162_out : STD_LOGIC;
	signal p163_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p163_out : STD_LOGIC;
	signal p164_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p164_out : STD_LOGIC;
	signal p165_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p165_out : STD_LOGIC;
	signal p166_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p166_out : STD_LOGIC;
	signal p167_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p167_out : STD_LOGIC;
	signal p168_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p168_out : STD_LOGIC;
	signal p169_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p169_out : STD_LOGIC;
	signal p170_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p170_out : STD_LOGIC;
	signal p171_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p171_out : STD_LOGIC;
	signal p172_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p172_out : STD_LOGIC;
	signal p173_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p173_out : STD_LOGIC;
	signal p174_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p174_out : STD_LOGIC;
	signal p175_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p175_out : STD_LOGIC;
	signal p176_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p176_out : STD_LOGIC;
	signal p177_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p177_out : STD_LOGIC;
	signal p178_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p178_out : STD_LOGIC;
	signal p179_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p179_out : STD_LOGIC;
	signal p180_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p180_out : STD_LOGIC;
	signal p181_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p181_out : STD_LOGIC;
	signal p182_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p182_out : STD_LOGIC;
	signal p183_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p183_out : STD_LOGIC;
	signal p184_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p184_out : STD_LOGIC;
	signal p185_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p185_out : STD_LOGIC;
	signal p186_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p186_out : STD_LOGIC;
	signal p187_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p187_out : STD_LOGIC;
	signal p188_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p188_out : STD_LOGIC;
	signal p189_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p189_out : STD_LOGIC;
	signal p190_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p190_out : STD_LOGIC;
	signal p191_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p191_out : STD_LOGIC;
	signal p192_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p192_out : STD_LOGIC;
	signal p193_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p193_out : STD_LOGIC;
	signal p194_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p194_out : STD_LOGIC;
	signal p195_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p195_out : STD_LOGIC;
	signal p196_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p196_out : STD_LOGIC;
	signal p197_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p197_out : STD_LOGIC;
	signal p198_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p198_out : STD_LOGIC;
	signal p199_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p199_out : STD_LOGIC;
	signal p200_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p200_out : STD_LOGIC;
	signal p201_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p201_out : STD_LOGIC;
	signal p202_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p202_out : STD_LOGIC;
	signal p203_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p203_out : STD_LOGIC;
	signal p204_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p204_out : STD_LOGIC;
	signal p205_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p205_out : STD_LOGIC;
	signal p206_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p206_out : STD_LOGIC;
	signal p207_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p207_out : STD_LOGIC;
	signal p208_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p208_out : STD_LOGIC;
	signal p209_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p209_out : STD_LOGIC;
	signal p210_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p210_out : STD_LOGIC;
	signal p211_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p211_out : STD_LOGIC;
	signal p212_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p212_out : STD_LOGIC;
	signal p213_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p213_out : STD_LOGIC;
	signal p214_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p214_out : STD_LOGIC;
	signal p215_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p215_out : STD_LOGIC;
	signal p216_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p216_out : STD_LOGIC;
	signal p217_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p217_out : STD_LOGIC;
	signal p218_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p218_out : STD_LOGIC;
	signal p219_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p219_out : STD_LOGIC;
	signal p220_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p220_out : STD_LOGIC;
	signal p221_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p221_out : STD_LOGIC;
	signal p222_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p222_out : STD_LOGIC;
	signal p223_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p223_out : STD_LOGIC;
	signal p224_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p224_out : STD_LOGIC;
	signal p225_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p225_out : STD_LOGIC;
	signal p226_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p226_out : STD_LOGIC;
	signal p227_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p227_out : STD_LOGIC;
	signal p228_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p228_out : STD_LOGIC;
	signal p229_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p229_out : STD_LOGIC;
	signal p230_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p230_out : STD_LOGIC;
	signal p231_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p231_out : STD_LOGIC;
	signal p232_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p232_out : STD_LOGIC;
	signal p233_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p233_out : STD_LOGIC;
	signal p234_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p234_out : STD_LOGIC;
	signal p235_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p235_out : STD_LOGIC;
	signal p236_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p236_out : STD_LOGIC;
	signal p237_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p237_out : STD_LOGIC;
	signal p238_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p238_out : STD_LOGIC;
	signal p239_in : STD_LOGIC_VECTOR(0 to 3 - 1);
	signal p239_out : STD_LOGIC;
	signal p240_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p240_out : STD_LOGIC;
	signal p241_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p241_out : STD_LOGIC;
	signal p242_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p242_out : STD_LOGIC;
	signal p243_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p243_out : STD_LOGIC;
	signal p244_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p244_out : STD_LOGIC;
	signal p245_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p245_out : STD_LOGIC;
	signal p246_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p246_out : STD_LOGIC;
	signal p247_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p247_out : STD_LOGIC;
	signal p248_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p248_out : STD_LOGIC;
	signal p249_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p249_out : STD_LOGIC;
	signal p250_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p250_out : STD_LOGIC;
	signal p251_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p251_out : STD_LOGIC;
	signal p252_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p252_out : STD_LOGIC;
	signal p253_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p253_out : STD_LOGIC;
	signal p254_in : STD_LOGIC_VECTOR(0 to 1 - 1);
	signal p254_out : STD_LOGIC;
	signal p255_in : STD_LOGIC_VECTOR(0 to 2 - 1);
	signal p255_out : STD_LOGIC;
	
    
    -- Dummies
    signal dummy0 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy1 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy2 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy3 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy4 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy5 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy6 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy7 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy8 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy9 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy10 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy11 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy12 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy13 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy14 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy15 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy16 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy17 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy18 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy19 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy20 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy21 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy22 : STD_LOGIC_VECTOR(0 to 11 - 2);
	signal dummy23 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy24 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy25 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy26 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy27 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy28 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy29 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy30 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy31 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy32 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy33 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy34 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy35 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy36 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy37 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy38 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy39 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy40 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy41 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy42 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy43 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy44 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy45 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy46 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy47 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy48 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy49 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy50 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy51 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy52 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy53 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy54 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy55 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy56 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy57 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy58 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy59 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy60 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy61 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy62 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy63 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy64 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy65 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy66 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy67 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy68 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy69 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy70 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy71 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy72 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy73 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy74 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy75 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy76 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy77 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy78 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy79 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy80 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy81 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy82 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy83 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy84 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy85 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy86 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy87 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy88 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy89 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy90 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy91 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy92 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy93 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy94 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy95 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy96 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy97 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy98 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy99 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy100 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy101 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy102 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy103 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy104 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy105 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy106 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy107 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy108 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy109 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy110 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy111 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy112 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy113 : STD_LOGIC_VECTOR(0 to 11 - 2);
	signal dummy114 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy115 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy116 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy117 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy118 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy119 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy120 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy121 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy122 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy123 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy124 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy125 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy126 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy127 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy128 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy129 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy130 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy131 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy132 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy133 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy134 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy135 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy136 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy137 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy138 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy139 : STD_LOGIC_VECTOR(0 to 11 - 2);
	signal dummy140 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy141 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy142 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy143 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy144 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy145 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy146 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy147 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy148 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy149 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy150 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy151 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy152 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy153 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy154 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy155 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy156 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy157 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy158 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy159 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy160 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy161 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy162 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy163 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy164 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy165 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy166 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy167 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy168 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy169 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy170 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy171 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy172 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy173 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy174 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy175 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy176 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy177 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy178 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy179 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy180 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy181 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy182 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy183 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy184 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy185 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy186 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy187 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy188 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy189 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy190 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy191 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy192 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy193 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy194 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy195 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy196 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy197 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy198 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy199 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy200 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy201 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy202 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy203 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy204 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy205 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy206 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy207 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy208 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy209 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy210 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy211 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy212 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy213 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy214 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy215 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy216 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy217 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy218 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy219 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy220 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy221 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy222 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy223 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy224 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy225 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy226 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy227 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy228 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy229 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy230 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy231 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy232 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy233 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy234 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy235 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy236 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy237 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy238 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy239 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy240 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy241 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy242 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy243 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy244 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy245 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy246 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy247 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy248 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy249 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy250 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy251 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy252 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy253 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy254 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy255 : STD_LOGIC_VECTOR(0 to 13 - 2);
	 

begin

    
    p0_in <= x(53) & x(80) & x(199);
    y(0) <= not(p0_out);
    p0 : perceptron
        Generic map (
            WEIGHTS => "100",
            SHIFT => 6,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p0_in,
            y(0) => p0_out,
            y(1 to 13 - 1) => dummy0
        );


    p1_in <= x(33) & x(80);
    y(1) <= not(p1_out);
    p1 : perceptron
        Generic map (
            WEIGHTS => "00",
            SHIFT => 6,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p1_in,
            y(0) => p1_out,
            y(1 to 12 - 1) => dummy1
        );


    p2_in(0) <= x(235);
    y(2) <= not(p2_out);
    p2 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => 9,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p2_in,
            y(0) => p2_out,
            y(1 to 12 - 1) => dummy2
        );


    p3_in(0) <= x(134);
    y(3) <= not(p3_out);
    p3 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p3_in,
            y(0) => p3_out,
            y(1 to 12 - 1) => dummy3
        );


    p4_in(0) <= x(134);
    y(4) <= not(p4_out);
    p4 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p4_in,
            y(0) => p4_out,
            y(1 to 12 - 1) => dummy4
        );


    p5_in(0) <= x(179);
    y(5) <= not(p5_out);
    p5 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => -36,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p5_in,
            y(0) => p5_out,
            y(1 to 12 - 1) => dummy5
        );


    p6_in(0) <= x(57);
    y(6) <= not(p6_out);
    p6 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p6_in,
            y(0) => p6_out,
            y(1 to 12 - 1) => dummy6
        );


    p7_in(0) <= x(80);
    y(7) <= not(p7_out);
    p7 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => 5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p7_in,
            y(0) => p7_out,
            y(1 to 12 - 1) => dummy7
        );


    p8_in(0) <= x(187);
    y(8) <= not(p8_out);
    p8 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => -10,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p8_in,
            y(0) => p8_out,
            y(1 to 12 - 1) => dummy8
        );


    p9_in <= x(26) & x(73) & x(189);
    y(9) <= not(p9_out);
    p9 : perceptron
        Generic map (
            WEIGHTS => "001",
            SHIFT => 6,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p9_in,
            y(0) => p9_out,
            y(1 to 13 - 1) => dummy9
        );


    p10_in <= x(53) & x(95);
    y(10) <= not(p10_out);
    p10 : perceptron
        Generic map (
            WEIGHTS => "11",
            SHIFT => 6,
            B => 7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p10_in,
            y(0) => p10_out,
            y(1 to 12 - 1) => dummy10
        );


    p11_in <= x(6) & x(9) & x(33) & x(117);
    y(11) <= not(p11_out);
    p11 : perceptron
        Generic map (
            WEIGHTS => "0011",
            SHIFT => 6,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p11_in,
            y(0) => p11_out,
            y(1 to 13 - 1) => dummy11
        );


    p12_in <= x(111) & x(239);
    y(12) <= not(p12_out);
    p12 : perceptron
        Generic map (
            WEIGHTS => "10",
            SHIFT => 7,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p12_in,
            y(0) => p12_out,
            y(1 to 13 - 1) => dummy12
        );


    p13_in(0) <= x(157);
    y(13) <= not(p13_out);
    p13 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => -10,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p13_in,
            y(0) => p13_out,
            y(1 to 12 - 1) => dummy13
        );


    p14_in(0) <= x(111);
    y(14) <= not(p14_out);
    p14 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p14_in,
            y(0) => p14_out,
            y(1 to 12 - 1) => dummy14
        );


    p15_in <= x(9) & x(50) & x(111) & x(182);
    y(15) <= not(p15_out);
    p15 : perceptron
        Generic map (
            WEIGHTS => "0010",
            SHIFT => 6,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p15_in,
            y(0) => p15_out,
            y(1 to 13 - 1) => dummy15
        );


    p16_in <= x(7) & x(45) & x(236) & x(251);
    y(16) <= not(p16_out);
    p16 : perceptron
        Generic map (
            WEIGHTS => "0001",
            SHIFT => 6,
            B => -7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p16_in,
            y(0) => p16_out,
            y(1 to 13 - 1) => dummy16
        );


    p17_in <= x(96) & x(143) & x(183) & x(195);
    y(17) <= not(p17_out);
    p17 : perceptron
        Generic map (
            WEIGHTS => "0011",
            SHIFT => 6,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p17_in,
            y(0) => p17_out,
            y(1 to 14 - 1) => dummy17
        );


    p18_in <= x(38) & x(126) & x(143);
    y(18) <= not(p18_out);
    p18 : perceptron
        Generic map (
            WEIGHTS => "000",
            SHIFT => 6,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p18_in,
            y(0) => p18_out,
            y(1 to 13 - 1) => dummy18
        );


    p19_in <= x(29) & x(128);
    y(19) <= not(p19_out);
    p19 : perceptron
        Generic map (
            WEIGHTS => "10",
            SHIFT => 6,
            B => -11,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p19_in,
            y(0) => p19_out,
            y(1 to 12 - 1) => dummy19
        );


    p20_in(0) <= x(40);
    y(20) <= not(p20_out);
    p20 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => 6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p20_in,
            y(0) => p20_out,
            y(1 to 12 - 1) => dummy20
        );


    p21_in(0) <= x(42);
    y(21) <= not(p21_out);
    p21 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => -13,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p21_in,
            y(0) => p21_out,
            y(1 to 12 - 1) => dummy21
        );


    p22_in(0) <= x(202);
    y(22) <= not(p22_out);
    p22 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 6,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p22_in,
            y(0) => p22_out,
            y(1 to 11 - 1) => dummy22
        );


    p23_in(0) <= x(61);
    y(23) <= not(p23_out);
    p23 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => 8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p23_in,
            y(0) => p23_out,
            y(1 to 12 - 1) => dummy23
        );


    p24_in <= x(40) & x(187) & x(228);
    y(24) <= not(p24_out);
    p24 : perceptron
        Generic map (
            WEIGHTS => "101",
            SHIFT => 6,
            B => 6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p24_in,
            y(0) => p24_out,
            y(1 to 13 - 1) => dummy24
        );


    p25_in <= x(9) & x(53) & x(91) & x(146);
    y(25) <= not(p25_out);
    p25 : perceptron
        Generic map (
            WEIGHTS => "1111",
            SHIFT => 6,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p25_in,
            y(0) => p25_out,
            y(1 to 13 - 1) => dummy25
        );


    p26_in(0) <= x(249);
    y(26) <= not(p26_out);
    p26 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => 9,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p26_in,
            y(0) => p26_out,
            y(1 to 12 - 1) => dummy26
        );


    p27_in <= x(80) & x(86) & x(164);
    y(27) <= not(p27_out);
    p27 : perceptron
        Generic map (
            WEIGHTS => "101",
            SHIFT => 6,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p27_in,
            y(0) => p27_out,
            y(1 to 13 - 1) => dummy27
        );


    p28_in(0) <= x(103);
    y(28) <= not(p28_out);
    p28 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => 11,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p28_in,
            y(0) => p28_out,
            y(1 to 12 - 1) => dummy28
        );


    p29_in <= x(50) & x(53) & x(60) & x(140) & x(204);
    y(29) <= not(p29_out);
    p29 : perceptron
        Generic map (
            WEIGHTS => "01000",
            SHIFT => 6,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p29_in,
            y(0) => p29_out,
            y(1 to 14 - 1) => dummy29
        );


    p30_in <= x(26) & x(130) & x(222);
    y(30) <= not(p30_out);
    p30 : perceptron
        Generic map (
            WEIGHTS => "111",
            SHIFT => 6,
            B => 4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p30_in,
            y(0) => p30_out,
            y(1 to 13 - 1) => dummy30
        );


    p31_in <= x(38) & x(66) & x(133) & x(204);
    y(31) <= not(p31_out);
    p31 : perceptron
        Generic map (
            WEIGHTS => "1101",
            SHIFT => 5,
            B => 4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p31_in,
            y(0) => p31_out,
            y(1 to 12 - 1) => dummy31
        );


    p32_in(0) <= x(191);
    y(32) <= not(p32_out);
    p32 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => 8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p32_in,
            y(0) => p32_out,
            y(1 to 12 - 1) => dummy32
        );


    p33_in <= x(126) & x(157);
    y(33) <= not(p33_out);
    p33 : perceptron
        Generic map (
            WEIGHTS => "11",
            SHIFT => 7,
            B => 4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p33_in,
            y(0) => p33_out,
            y(1 to 13 - 1) => dummy33
        );


    p34_in <= x(9) & x(53) & x(65);
    y(34) <= not(p34_out);
    p34 : perceptron
        Generic map (
            WEIGHTS => "011",
            SHIFT => 6,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p34_in,
            y(0) => p34_out,
            y(1 to 13 - 1) => dummy34
        );


    p35_in(0) <= x(107);
    y(35) <= not(p35_out);
    p35 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => 5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p35_in,
            y(0) => p35_out,
            y(1 to 12 - 1) => dummy35
        );


    p36_in <= x(7) & x(45);
    y(36) <= not(p36_out);
    p36 : perceptron
        Generic map (
            WEIGHTS => "00",
            SHIFT => 7,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p36_in,
            y(0) => p36_out,
            y(1 to 13 - 1) => dummy36
        );


    p37_in <= x(86) & x(227) & x(236);
    y(37) <= not(p37_out);
    p37 : perceptron
        Generic map (
            WEIGHTS => "010",
            SHIFT => 6,
            B => -10,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p37_in,
            y(0) => p37_out,
            y(1 to 13 - 1) => dummy37
        );


    p38_in <= x(13) & x(45) & x(101) & x(162);
    y(38) <= not(p38_out);
    p38 : perceptron
        Generic map (
            WEIGHTS => "1011",
            SHIFT => 6,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p38_in,
            y(0) => p38_out,
            y(1 to 13 - 1) => dummy38
        );


    p39_in(0) <= x(192);
    y(39) <= not(p39_out);
    p39 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => 14,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p39_in,
            y(0) => p39_out,
            y(1 to 12 - 1) => dummy39
        );


    p40_in <= x(117) & x(189) & x(249);
    y(40) <= not(p40_out);
    p40 : perceptron
        Generic map (
            WEIGHTS => "010",
            SHIFT => 6,
            B => 8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p40_in,
            y(0) => p40_out,
            y(1 to 13 - 1) => dummy40
        );


    p41_in <= x(8) & x(202);
    y(41) <= not(p41_out);
    p41 : perceptron
        Generic map (
            WEIGHTS => "00",
            SHIFT => 6,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p41_in,
            y(0) => p41_out,
            y(1 to 12 - 1) => dummy41
        );


    p42_in <= x(31) & x(239);
    y(42) <= not(p42_out);
    p42 : perceptron
        Generic map (
            WEIGHTS => "00",
            SHIFT => 6,
            B => -8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p42_in,
            y(0) => p42_out,
            y(1 to 12 - 1) => dummy42
        );


    p43_in <= x(56) & x(184) & x(226);
    y(43) <= not(p43_out);
    p43 : perceptron
        Generic map (
            WEIGHTS => "111",
            SHIFT => 6,
            B => 7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p43_in,
            y(0) => p43_out,
            y(1 to 13 - 1) => dummy43
        );


    p44_in(0) <= x(130);
    y(44) <= not(p44_out);
    p44 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p44_in,
            y(0) => p44_out,
            y(1 to 12 - 1) => dummy44
        );


    p45_in(0) <= x(198);
    y(45) <= not(p45_out);
    p45 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => 12,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p45_in,
            y(0) => p45_out,
            y(1 to 12 - 1) => dummy45
        );


    p46_in <= x(92) & x(130) & x(211) & x(244);
    y(46) <= not(p46_out);
    p46 : perceptron
        Generic map (
            WEIGHTS => "1100",
            SHIFT => 6,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p46_in,
            y(0) => p46_out,
            y(1 to 14 - 1) => dummy46
        );


    p47_in(0) <= x(32);
    y(47) <= not(p47_out);
    p47 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p47_in,
            y(0) => p47_out,
            y(1 to 12 - 1) => dummy47
        );


    p48_in(0) <= x(111);
    y(48) <= not(p48_out);
    p48 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p48_in,
            y(0) => p48_out,
            y(1 to 12 - 1) => dummy48
        );


    p49_in(0) <= x(60);
    y(49) <= not(p49_out);
    p49 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p49_in,
            y(0) => p49_out,
            y(1 to 12 - 1) => dummy49
        );


    p50_in(0) <= x(95);
    y(50) <= not(p50_out);
    p50 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => 12,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p50_in,
            y(0) => p50_out,
            y(1 to 12 - 1) => dummy50
        );


    p51_in <= x(7) & x(115) & x(143);
    y(51) <= not(p51_out);
    p51 : perceptron
        Generic map (
            WEIGHTS => "110",
            SHIFT => 6,
            B => 19,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p51_in,
            y(0) => p51_out,
            y(1 to 13 - 1) => dummy51
        );


    p52_in(0) <= x(48);
    y(52) <= not(p52_out);
    p52 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p52_in,
            y(0) => p52_out,
            y(1 to 12 - 1) => dummy52
        );


    p53_in <= x(80) & x(168) & x(250);
    y(53) <= not(p53_out);
    p53 : perceptron
        Generic map (
            WEIGHTS => "110",
            SHIFT => 6,
            B => 4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p53_in,
            y(0) => p53_out,
            y(1 to 13 - 1) => dummy53
        );


    p54_in <= x(53) & x(129) & x(212);
    y(54) <= not(p54_out);
    p54 : perceptron
        Generic map (
            WEIGHTS => "000",
            SHIFT => 6,
            B => 13,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p54_in,
            y(0) => p54_out,
            y(1 to 13 - 1) => dummy54
        );


    p55_in(0) <= x(103);
    y(55) <= not(p55_out);
    p55 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => 11,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p55_in,
            y(0) => p55_out,
            y(1 to 12 - 1) => dummy55
        );


    p56_in <= x(47) & x(73);
    y(56) <= not(p56_out);
    p56 : perceptron
        Generic map (
            WEIGHTS => "10",
            SHIFT => 6,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p56_in,
            y(0) => p56_out,
            y(1 to 12 - 1) => dummy56
        );


    p57_in <= x(32) & x(53) & x(158);
    y(57) <= not(p57_out);
    p57 : perceptron
        Generic map (
            WEIGHTS => "010",
            SHIFT => 6,
            B => 4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p57_in,
            y(0) => p57_out,
            y(1 to 13 - 1) => dummy57
        );


    p58_in <= x(80) & x(160) & x(162);
    y(58) <= not(p58_out);
    p58 : perceptron
        Generic map (
            WEIGHTS => "011",
            SHIFT => 6,
            B => -8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p58_in,
            y(0) => p58_out,
            y(1 to 13 - 1) => dummy58
        );


    p59_in(0) <= x(229);
    y(59) <= not(p59_out);
    p59 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => 8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p59_in,
            y(0) => p59_out,
            y(1 to 12 - 1) => dummy59
        );


    p60_in <= x(6) & x(95);
    y(60) <= not(p60_out);
    p60 : perceptron
        Generic map (
            WEIGHTS => "01",
            SHIFT => 6,
            B => 10,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p60_in,
            y(0) => p60_out,
            y(1 to 12 - 1) => dummy60
        );


    p61_in <= x(33) & x(59) & x(86) & x(96) & x(184) & x(216);
    y(61) <= not(p61_out);
    p61 : perceptron
        Generic map (
            WEIGHTS => "101001",
            SHIFT => 5,
            B => -14,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p61_in,
            y(0) => p61_out,
            y(1 to 13 - 1) => dummy61
        );


    p62_in <= x(61) & x(80) & x(227) & x(236);
    y(62) <= not(p62_out);
    p62 : perceptron
        Generic map (
            WEIGHTS => "1101",
            SHIFT => 6,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p62_in,
            y(0) => p62_out,
            y(1 to 13 - 1) => dummy62
        );


    p63_in <= x(56) & x(130) & x(226);
    y(63) <= not(p63_out);
    p63 : perceptron
        Generic map (
            WEIGHTS => "101",
            SHIFT => 6,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p63_in,
            y(0) => p63_out,
            y(1 to 13 - 1) => dummy63
        );


    p64_in(0) <= x(184);
    y(64) <= not(p64_out);
    p64 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => 6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p64_in,
            y(0) => p64_out,
            y(1 to 12 - 1) => dummy64
        );


    p65_in(0) <= x(111);
    y(65) <= not(p65_out);
    p65 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p65_in,
            y(0) => p65_out,
            y(1 to 12 - 1) => dummy65
        );


    p66_in <= x(88) & x(195) & x(217);
    y(66) <= not(p66_out);
    p66 : perceptron
        Generic map (
            WEIGHTS => "011",
            SHIFT => 6,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p66_in,
            y(0) => p66_out,
            y(1 to 13 - 1) => dummy66
        );


    p67_in <= x(126) & x(143) & x(191);
    y(67) <= not(p67_out);
    p67 : perceptron
        Generic map (
            WEIGHTS => "000",
            SHIFT => 6,
            B => -6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p67_in,
            y(0) => p67_out,
            y(1 to 13 - 1) => dummy67
        );


    p68_in <= x(119) & x(177) & x(234);
    y(68) <= not(p68_out);
    p68 : perceptron
        Generic map (
            WEIGHTS => "000",
            SHIFT => 6,
            B => -6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p68_in,
            y(0) => p68_out,
            y(1 to 13 - 1) => dummy68
        );


    p69_in <= x(45) & x(228);
    y(69) <= not(p69_out);
    p69 : perceptron
        Generic map (
            WEIGHTS => "01",
            SHIFT => 6,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p69_in,
            y(0) => p69_out,
            y(1 to 12 - 1) => dummy69
        );


    p70_in <= x(30) & x(105) & x(237);
    y(70) <= not(p70_out);
    p70 : perceptron
        Generic map (
            WEIGHTS => "101",
            SHIFT => 6,
            B => 8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p70_in,
            y(0) => p70_out,
            y(1 to 13 - 1) => dummy70
        );


    p71_in <= x(59) & x(144);
    y(71) <= not(p71_out);
    p71 : perceptron
        Generic map (
            WEIGHTS => "10",
            SHIFT => 6,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p71_in,
            y(0) => p71_out,
            y(1 to 12 - 1) => dummy71
        );


    p72_in <= x(60) & x(197);
    y(72) <= not(p72_out);
    p72 : perceptron
        Generic map (
            WEIGHTS => "01",
            SHIFT => 6,
            B => -12,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p72_in,
            y(0) => p72_out,
            y(1 to 12 - 1) => dummy72
        );


    p73_in <= x(62) & x(75) & x(80);
    y(73) <= not(p73_out);
    p73 : perceptron
        Generic map (
            WEIGHTS => "111",
            SHIFT => 6,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p73_in,
            y(0) => p73_out,
            y(1 to 13 - 1) => dummy73
        );


    p74_in <= x(22) & x(160) & x(162);
    y(74) <= not(p74_out);
    p74 : perceptron
        Generic map (
            WEIGHTS => "011",
            SHIFT => 6,
            B => -14,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p74_in,
            y(0) => p74_out,
            y(1 to 13 - 1) => dummy74
        );


    p75_in(0) <= x(125);
    y(75) <= not(p75_out);
    p75 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => 13,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p75_in,
            y(0) => p75_out,
            y(1 to 12 - 1) => dummy75
        );


    p76_in(0) <= x(193);
    y(76) <= not(p76_out);
    p76 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => 12,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p76_in,
            y(0) => p76_out,
            y(1 to 12 - 1) => dummy76
        );


    p77_in <= x(86) & x(184);
    y(77) <= not(p77_out);
    p77 : perceptron
        Generic map (
            WEIGHTS => "10",
            SHIFT => 6,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p77_in,
            y(0) => p77_out,
            y(1 to 12 - 1) => dummy77
        );


    p78_in <= x(78) & x(166) & x(184);
    y(78) <= not(p78_out);
    p78 : perceptron
        Generic map (
            WEIGHTS => "011",
            SHIFT => 6,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p78_in,
            y(0) => p78_out,
            y(1 to 13 - 1) => dummy78
        );


    p79_in <= x(153) & x(198);
    y(79) <= not(p79_out);
    p79 : perceptron
        Generic map (
            WEIGHTS => "11",
            SHIFT => 6,
            B => -8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p79_in,
            y(0) => p79_out,
            y(1 to 12 - 1) => dummy79
        );


    p80_in(0) <= x(22);
    y(80) <= not(p80_out);
    p80 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => 13,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p80_in,
            y(0) => p80_out,
            y(1 to 12 - 1) => dummy80
        );


    p81_in(0) <= x(160);
    y(81) <= not(p81_out);
    p81 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => -21,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p81_in,
            y(0) => p81_out,
            y(1 to 12 - 1) => dummy81
        );


    p82_in(0) <= x(103);
    y(82) <= not(p82_out);
    p82 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => 11,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p82_in,
            y(0) => p82_out,
            y(1 to 12 - 1) => dummy82
        );


    p83_in <= x(86) & x(112) & x(183);
    y(83) <= not(p83_out);
    p83 : perceptron
        Generic map (
            WEIGHTS => "111",
            SHIFT => 6,
            B => 13,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p83_in,
            y(0) => p83_out,
            y(1 to 13 - 1) => dummy83
        );


    p84_in <= x(7) & x(45) & x(216) & x(230) & x(236);
    y(84) <= not(p84_out);
    p84 : perceptron
        Generic map (
            WEIGHTS => "00000",
            SHIFT => 6,
            B => -6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p84_in,
            y(0) => p84_out,
            y(1 to 14 - 1) => dummy84
        );


    p85_in <= x(50) & x(92) & x(214) & x(244);
    y(85) <= not(p85_out);
    p85 : perceptron
        Generic map (
            WEIGHTS => "1100",
            SHIFT => 6,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p85_in,
            y(0) => p85_out,
            y(1 to 13 - 1) => dummy85
        );


    p86_in <= x(22) & x(133) & x(184);
    y(86) <= not(p86_out);
    p86 : perceptron
        Generic map (
            WEIGHTS => "110",
            SHIFT => 6,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p86_in,
            y(0) => p86_out,
            y(1 to 13 - 1) => dummy86
        );


    p87_in <= x(80) & x(91);
    y(87) <= not(p87_out);
    p87 : perceptron
        Generic map (
            WEIGHTS => "00",
            SHIFT => 6,
            B => -6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p87_in,
            y(0) => p87_out,
            y(1 to 12 - 1) => dummy87
        );


    p88_in <= x(19) & x(129) & x(137);
    y(88) <= not(p88_out);
    p88 : perceptron
        Generic map (
            WEIGHTS => "100",
            SHIFT => 6,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p88_in,
            y(0) => p88_out,
            y(1 to 13 - 1) => dummy88
        );


    p89_in <= x(45) & x(137);
    y(89) <= not(p89_out);
    p89 : perceptron
        Generic map (
            WEIGHTS => "11",
            SHIFT => 6,
            B => 6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p89_in,
            y(0) => p89_out,
            y(1 to 12 - 1) => dummy89
        );


    p90_in(0) <= x(13);
    y(90) <= not(p90_out);
    p90 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => -9,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p90_in,
            y(0) => p90_out,
            y(1 to 12 - 1) => dummy90
        );


    p91_in(0) <= x(235);
    y(91) <= not(p91_out);
    p91 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => 13,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p91_in,
            y(0) => p91_out,
            y(1 to 12 - 1) => dummy91
        );


    p92_in <= x(27) & x(33) & x(140);
    y(92) <= not(p92_out);
    p92 : perceptron
        Generic map (
            WEIGHTS => "101",
            SHIFT => 6,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p92_in,
            y(0) => p92_out,
            y(1 to 13 - 1) => dummy92
        );


    p93_in(0) <= x(103);
    y(93) <= not(p93_out);
    p93 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => 11,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p93_in,
            y(0) => p93_out,
            y(1 to 12 - 1) => dummy93
        );


    p94_in <= x(38) & x(101) & x(239);
    y(94) <= not(p94_out);
    p94 : perceptron
        Generic map (
            WEIGHTS => "100",
            SHIFT => 6,
            B => 6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p94_in,
            y(0) => p94_out,
            y(1 to 13 - 1) => dummy94
        );


    p95_in <= x(19) & x(91) & x(205);
    y(95) <= not(p95_out);
    p95 : perceptron
        Generic map (
            WEIGHTS => "011",
            SHIFT => 6,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p95_in,
            y(0) => p95_out,
            y(1 to 13 - 1) => dummy95
        );


    p96_in <= x(9) & x(113) & x(235);
    y(96) <= not(p96_out);
    p96 : perceptron
        Generic map (
            WEIGHTS => "001",
            SHIFT => 6,
            B => -14,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p96_in,
            y(0) => p96_out,
            y(1 to 13 - 1) => dummy96
        );


    p97_in <= x(150) & x(203);
    y(97) <= not(p97_out);
    p97 : perceptron
        Generic map (
            WEIGHTS => "00",
            SHIFT => 6,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p97_in,
            y(0) => p97_out,
            y(1 to 12 - 1) => dummy97
        );


    p98_in <= x(8) & x(39);
    y(98) <= not(p98_out);
    p98 : perceptron
        Generic map (
            WEIGHTS => "01",
            SHIFT => 6,
            B => 15,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p98_in,
            y(0) => p98_out,
            y(1 to 12 - 1) => dummy98
        );


    p99_in <= x(117) & x(119);
    y(99) <= not(p99_out);
    p99 : perceptron
        Generic map (
            WEIGHTS => "01",
            SHIFT => 6,
            B => 6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p99_in,
            y(0) => p99_out,
            y(1 to 12 - 1) => dummy99
        );


    p100_in(0) <= x(192);
    y(100) <= not(p100_out);
    p100 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => -15,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p100_in,
            y(0) => p100_out,
            y(1 to 12 - 1) => dummy100
        );


    p101_in <= x(137) & x(222);
    y(101) <= not(p101_out);
    p101 : perceptron
        Generic map (
            WEIGHTS => "00",
            SHIFT => 6,
            B => -8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p101_in,
            y(0) => p101_out,
            y(1 to 12 - 1) => dummy101
        );


    p102_in <= x(19) & x(143);
    y(102) <= not(p102_out);
    p102 : perceptron
        Generic map (
            WEIGHTS => "01",
            SHIFT => 6,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p102_in,
            y(0) => p102_out,
            y(1 to 12 - 1) => dummy102
        );


    p103_in <= x(76) & x(163);
    y(103) <= not(p103_out);
    p103 : perceptron
        Generic map (
            WEIGHTS => "00",
            SHIFT => 6,
            B => 4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p103_in,
            y(0) => p103_out,
            y(1 to 12 - 1) => dummy103
        );


    p104_in <= x(8) & x(33);
    y(104) <= not(p104_out);
    p104 : perceptron
        Generic map (
            WEIGHTS => "01",
            SHIFT => 7,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p104_in,
            y(0) => p104_out,
            y(1 to 13 - 1) => dummy104
        );


    p105_in <= x(13) & x(22) & x(100) & x(228);
    y(105) <= not(p105_out);
    p105 : perceptron
        Generic map (
            WEIGHTS => "0010",
            SHIFT => 5,
            B => -10,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p105_in,
            y(0) => p105_out,
            y(1 to 12 - 1) => dummy105
        );


    p106_in <= x(82) & x(130);
    y(106) <= not(p106_out);
    p106 : perceptron
        Generic map (
            WEIGHTS => "00",
            SHIFT => 6,
            B => -13,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p106_in,
            y(0) => p106_out,
            y(1 to 12 - 1) => dummy106
        );


    p107_in(0) <= x(132);
    y(107) <= not(p107_out);
    p107 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p107_in,
            y(0) => p107_out,
            y(1 to 12 - 1) => dummy107
        );


    p108_in(0) <= x(172);
    y(108) <= not(p108_out);
    p108 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => -15,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p108_in,
            y(0) => p108_out,
            y(1 to 12 - 1) => dummy108
        );


    p109_in <= x(39) & x(203) & x(204) & x(239);
    y(109) <= not(p109_out);
    p109 : perceptron
        Generic map (
            WEIGHTS => "1110",
            SHIFT => 6,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p109_in,
            y(0) => p109_out,
            y(1 to 14 - 1) => dummy109
        );


    p110_in(0) <= x(193);
    y(110) <= not(p110_out);
    p110 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => -13,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p110_in,
            y(0) => p110_out,
            y(1 to 12 - 1) => dummy110
        );


    p111_in <= x(105) & x(249);
    y(111) <= not(p111_out);
    p111 : perceptron
        Generic map (
            WEIGHTS => "01",
            SHIFT => 7,
            B => -9,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p111_in,
            y(0) => p111_out,
            y(1 to 13 - 1) => dummy111
        );


    p112_in <= x(45) & x(122) & x(213);
    y(112) <= not(p112_out);
    p112 : perceptron
        Generic map (
            WEIGHTS => "101",
            SHIFT => 6,
            B => 5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p112_in,
            y(0) => p112_out,
            y(1 to 13 - 1) => dummy112
        );


    p113_in(0) <= x(30);
    y(113) <= not(p113_out);
    p113 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 6,
            B => 11,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p113_in,
            y(0) => p113_out,
            y(1 to 11 - 1) => dummy113
        );


    p114_in <= x(29) & x(89) & x(194);
    y(114) <= not(p114_out);
    p114 : perceptron
        Generic map (
            WEIGHTS => "010",
            SHIFT => 6,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p114_in,
            y(0) => p114_out,
            y(1 to 13 - 1) => dummy114
        );


    p115_in(0) <= x(105);
    y(115) <= not(p115_out);
    p115 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p115_in,
            y(0) => p115_out,
            y(1 to 12 - 1) => dummy115
        );


    p116_in(0) <= x(177);
    y(116) <= not(p116_out);
    p116 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p116_in,
            y(0) => p116_out,
            y(1 to 12 - 1) => dummy116
        );


    p117_in(0) <= x(177);
    y(117) <= not(p117_out);
    p117 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => 4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p117_in,
            y(0) => p117_out,
            y(1 to 12 - 1) => dummy117
        );


    p118_in(0) <= x(113);
    y(118) <= not(p118_out);
    p118 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => 9,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p118_in,
            y(0) => p118_out,
            y(1 to 12 - 1) => dummy118
        );


    p119_in(0) <= x(182);
    y(119) <= not(p119_out);
    p119 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => 5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p119_in,
            y(0) => p119_out,
            y(1 to 12 - 1) => dummy119
        );


    p120_in(0) <= x(184);
    y(120) <= not(p120_out);
    p120 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => -7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p120_in,
            y(0) => p120_out,
            y(1 to 12 - 1) => dummy120
        );


    p121_in <= x(19) & x(143);
    y(121) <= not(p121_out);
    p121 : perceptron
        Generic map (
            WEIGHTS => "01",
            SHIFT => 6,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p121_in,
            y(0) => p121_out,
            y(1 to 12 - 1) => dummy121
        );


    p122_in <= x(15) & x(22) & x(130);
    y(122) <= not(p122_out);
    p122 : perceptron
        Generic map (
            WEIGHTS => "101",
            SHIFT => 6,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p122_in,
            y(0) => p122_out,
            y(1 to 13 - 1) => dummy122
        );


    p123_in(0) <= x(190);
    y(123) <= not(p123_out);
    p123 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => 10,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p123_in,
            y(0) => p123_out,
            y(1 to 12 - 1) => dummy123
        );


    p124_in <= x(62) & x(103);
    y(124) <= not(p124_out);
    p124 : perceptron
        Generic map (
            WEIGHTS => "10",
            SHIFT => 7,
            B => 12,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p124_in,
            y(0) => p124_out,
            y(1 to 13 - 1) => dummy124
        );


    p125_in <= x(59) & x(144);
    y(125) <= not(p125_out);
    p125 : perceptron
        Generic map (
            WEIGHTS => "10",
            SHIFT => 6,
            B => 4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p125_in,
            y(0) => p125_out,
            y(1 to 12 - 1) => dummy125
        );


    p126_in <= x(42) & x(175);
    y(126) <= not(p126_out);
    p126 : perceptron
        Generic map (
            WEIGHTS => "01",
            SHIFT => 6,
            B => -11,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p126_in,
            y(0) => p126_out,
            y(1 to 12 - 1) => dummy126
        );


    p127_in(0) <= x(239);
    y(127) <= not(p127_out);
    p127 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p127_in,
            y(0) => p127_out,
            y(1 to 12 - 1) => dummy127
        );


    p128_in(0) <= x(38);
    y(128) <= not(p128_out);
    p128 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p128_in,
            y(0) => p128_out,
            y(1 to 12 - 1) => dummy128
        );


    p129_in(0) <= x(196);
    y(129) <= not(p129_out);
    p129 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => -18,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p129_in,
            y(0) => p129_out,
            y(1 to 12 - 1) => dummy129
        );


    p130_in <= x(22) & x(197) & x(211) & x(229);
    y(130) <= not(p130_out);
    p130 : perceptron
        Generic map (
            WEIGHTS => "0011",
            SHIFT => 5,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p130_in,
            y(0) => p130_out,
            y(1 to 13 - 1) => dummy130
        );


    p131_in(0) <= x(239);
    y(131) <= not(p131_out);
    p131 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p131_in,
            y(0) => p131_out,
            y(1 to 12 - 1) => dummy131
        );


    p132_in <= x(50) & x(143) & x(229);
    y(132) <= not(p132_out);
    p132 : perceptron
        Generic map (
            WEIGHTS => "101",
            SHIFT => 6,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p132_in,
            y(0) => p132_out,
            y(1 to 13 - 1) => dummy132
        );


    p133_in <= x(75) & x(80) & x(204) & x(235);
    y(133) <= not(p133_out);
    p133 : perceptron
        Generic map (
            WEIGHTS => "0001",
            SHIFT => 6,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p133_in,
            y(0) => p133_out,
            y(1 to 13 - 1) => dummy133
        );


    p134_in <= x(33) & x(133);
    y(134) <= not(p134_out);
    p134 : perceptron
        Generic map (
            WEIGHTS => "00",
            SHIFT => 6,
            B => 5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p134_in,
            y(0) => p134_out,
            y(1 to 12 - 1) => dummy134
        );


    p135_in(0) <= x(42);
    y(135) <= not(p135_out);
    p135 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => 12,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p135_in,
            y(0) => p135_out,
            y(1 to 12 - 1) => dummy135
        );


    p136_in(0) <= x(134);
    y(136) <= not(p136_out);
    p136 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p136_in,
            y(0) => p136_out,
            y(1 to 12 - 1) => dummy136
        );


    p137_in(0) <= x(59);
    y(137) <= not(p137_out);
    p137 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p137_in,
            y(0) => p137_out,
            y(1 to 12 - 1) => dummy137
        );


    p138_in <= x(103) & x(171) & x(177) & x(240);
    y(138) <= not(p138_out);
    p138 : perceptron
        Generic map (
            WEIGHTS => "0010",
            SHIFT => 6,
            B => 7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p138_in,
            y(0) => p138_out,
            y(1 to 14 - 1) => dummy138
        );


    p139_in(0) <= x(56);
    y(139) <= not(p139_out);
    p139 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 6,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p139_in,
            y(0) => p139_out,
            y(1 to 11 - 1) => dummy139
        );


    p140_in <= x(118) & x(126);
    y(140) <= not(p140_out);
    p140 : perceptron
        Generic map (
            WEIGHTS => "01",
            SHIFT => 6,
            B => -11,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p140_in,
            y(0) => p140_out,
            y(1 to 12 - 1) => dummy140
        );


    p141_in <= x(189) & x(253);
    y(141) <= not(p141_out);
    p141 : perceptron
        Generic map (
            WEIGHTS => "01",
            SHIFT => 7,
            B => -7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p141_in,
            y(0) => p141_out,
            y(1 to 13 - 1) => dummy141
        );


    p142_in <= x(20) & x(250);
    y(142) <= not(p142_out);
    p142 : perceptron
        Generic map (
            WEIGHTS => "10",
            SHIFT => 6,
            B => 7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p142_in,
            y(0) => p142_out,
            y(1 to 12 - 1) => dummy142
        );


    p143_in <= x(60) & x(162);
    y(143) <= not(p143_out);
    p143 : perceptron
        Generic map (
            WEIGHTS => "00",
            SHIFT => 6,
            B => -6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p143_in,
            y(0) => p143_out,
            y(1 to 12 - 1) => dummy143
        );


    p144_in <= x(6) & x(103);
    y(144) <= not(p144_out);
    p144 : perceptron
        Generic map (
            WEIGHTS => "01",
            SHIFT => 7,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p144_in,
            y(0) => p144_out,
            y(1 to 13 - 1) => dummy144
        );


    p145_in <= x(19) & x(38);
    y(145) <= not(p145_out);
    p145 : perceptron
        Generic map (
            WEIGHTS => "01",
            SHIFT => 6,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p145_in,
            y(0) => p145_out,
            y(1 to 12 - 1) => dummy145
        );


    p146_in(0) <= x(13);
    y(146) <= not(p146_out);
    p146 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => 8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p146_in,
            y(0) => p146_out,
            y(1 to 12 - 1) => dummy146
        );


    p147_in(0) <= x(226);
    y(147) <= not(p147_out);
    p147 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p147_in,
            y(0) => p147_out,
            y(1 to 12 - 1) => dummy147
        );


    p148_in <= x(205) & x(217);
    y(148) <= not(p148_out);
    p148 : perceptron
        Generic map (
            WEIGHTS => "10",
            SHIFT => 6,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p148_in,
            y(0) => p148_out,
            y(1 to 12 - 1) => dummy148
        );


    p149_in <= x(19) & x(133) & x(184);
    y(149) <= not(p149_out);
    p149 : perceptron
        Generic map (
            WEIGHTS => "001",
            SHIFT => 6,
            B => 5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p149_in,
            y(0) => p149_out,
            y(1 to 13 - 1) => dummy149
        );


    p150_in(0) <= x(130);
    y(150) <= not(p150_out);
    p150 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => 4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p150_in,
            y(0) => p150_out,
            y(1 to 12 - 1) => dummy150
        );


    p151_in(0) <= x(253);
    y(151) <= not(p151_out);
    p151 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => 4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p151_in,
            y(0) => p151_out,
            y(1 to 12 - 1) => dummy151
        );


    p152_in(0) <= x(80);
    y(152) <= not(p152_out);
    p152 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => 5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p152_in,
            y(0) => p152_out,
            y(1 to 12 - 1) => dummy152
        );


    p153_in <= x(7) & x(91);
    y(153) <= not(p153_out);
    p153 : perceptron
        Generic map (
            WEIGHTS => "00",
            SHIFT => 6,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p153_in,
            y(0) => p153_out,
            y(1 to 12 - 1) => dummy153
        );


    p154_in(0) <= x(250);
    y(154) <= not(p154_out);
    p154 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p154_in,
            y(0) => p154_out,
            y(1 to 12 - 1) => dummy154
        );


    p155_in <= x(62) & x(103) & x(243);
    y(155) <= not(p155_out);
    p155 : perceptron
        Generic map (
            WEIGHTS => "011",
            SHIFT => 6,
            B => -9,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p155_in,
            y(0) => p155_out,
            y(1 to 13 - 1) => dummy155
        );


    p156_in <= x(7) & x(8) & x(38) & x(194);
    y(156) <= not(p156_out);
    p156 : perceptron
        Generic map (
            WEIGHTS => "1010",
            SHIFT => 5,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p156_in,
            y(0) => p156_out,
            y(1 to 12 - 1) => dummy156
        );


    p157_in(0) <= x(107);
    y(157) <= not(p157_out);
    p157 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => -6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p157_in,
            y(0) => p157_out,
            y(1 to 12 - 1) => dummy157
        );


    p158_in <= x(140) & x(184);
    y(158) <= not(p158_out);
    p158 : perceptron
        Generic map (
            WEIGHTS => "10",
            SHIFT => 6,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p158_in,
            y(0) => p158_out,
            y(1 to 12 - 1) => dummy158
        );


    p159_in <= x(81) & x(195) & x(204);
    y(159) <= not(p159_out);
    p159 : perceptron
        Generic map (
            WEIGHTS => "001",
            SHIFT => 6,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p159_in,
            y(0) => p159_out,
            y(1 to 13 - 1) => dummy159
        );


    p160_in <= x(81) & x(228);
    y(160) <= not(p160_out);
    p160 : perceptron
        Generic map (
            WEIGHTS => "10",
            SHIFT => 7,
            B => 7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p160_in,
            y(0) => p160_out,
            y(1 to 13 - 1) => dummy160
        );


    p161_in(0) <= x(79);
    y(161) <= not(p161_out);
    p161 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => 8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p161_in,
            y(0) => p161_out,
            y(1 to 12 - 1) => dummy161
        );


    p162_in(0) <= x(39);
    y(162) <= not(p162_out);
    p162 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => 22,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p162_in,
            y(0) => p162_out,
            y(1 to 12 - 1) => dummy162
        );


    p163_in(0) <= x(162);
    y(163) <= not(p163_out);
    p163 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => 6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p163_in,
            y(0) => p163_out,
            y(1 to 12 - 1) => dummy163
        );


    p164_in <= x(33) & x(91) & x(162);
    y(164) <= not(p164_out);
    p164 : perceptron
        Generic map (
            WEIGHTS => "111",
            SHIFT => 6,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p164_in,
            y(0) => p164_out,
            y(1 to 13 - 1) => dummy164
        );


    p165_in <= x(153) & x(189) & x(198);
    y(165) <= not(p165_out);
    p165 : perceptron
        Generic map (
            WEIGHTS => "101",
            SHIFT => 6,
            B => -8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p165_in,
            y(0) => p165_out,
            y(1 to 13 - 1) => dummy165
        );


    p166_in(0) <= x(249);
    y(166) <= not(p166_out);
    p166 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => 9,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p166_in,
            y(0) => p166_out,
            y(1 to 12 - 1) => dummy166
        );


    p167_in <= x(30) & x(73) & x(78) & x(153) & x(157);
    y(167) <= not(p167_out);
    p167 : perceptron
        Generic map (
            WEIGHTS => "10001",
            SHIFT => 6,
            B => 8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p167_in,
            y(0) => p167_out,
            y(1 to 14 - 1) => dummy167
        );


    p168_in <= x(33) & x(110) & x(247);
    y(168) <= not(p168_out);
    p168 : perceptron
        Generic map (
            WEIGHTS => "001",
            SHIFT => 6,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p168_in,
            y(0) => p168_out,
            y(1 to 13 - 1) => dummy168
        );


    p169_in <= x(50) & x(177);
    y(169) <= not(p169_out);
    p169 : perceptron
        Generic map (
            WEIGHTS => "10",
            SHIFT => 7,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p169_in,
            y(0) => p169_out,
            y(1 to 13 - 1) => dummy169
        );


    p170_in <= x(44) & x(164);
    y(170) <= not(p170_out);
    p170 : perceptron
        Generic map (
            WEIGHTS => "01",
            SHIFT => 6,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p170_in,
            y(0) => p170_out,
            y(1 to 12 - 1) => dummy170
        );


    p171_in <= x(96) & x(195);
    y(171) <= not(p171_out);
    p171 : perceptron
        Generic map (
            WEIGHTS => "10",
            SHIFT => 6,
            B => 11,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p171_in,
            y(0) => p171_out,
            y(1 to 12 - 1) => dummy171
        );


    p172_in <= x(184) & x(250);
    y(172) <= not(p172_out);
    p172 : perceptron
        Generic map (
            WEIGHTS => "10",
            SHIFT => 7,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p172_in,
            y(0) => p172_out,
            y(1 to 13 - 1) => dummy172
        );


    p173_in <= x(39) & x(97) & x(111) & x(143) & x(191);
    y(173) <= not(p173_out);
    p173 : perceptron
        Generic map (
            WEIGHTS => "00011",
            SHIFT => 5,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p173_in,
            y(0) => p173_out,
            y(1 to 13 - 1) => dummy173
        );


    p174_in <= x(119) & x(143);
    y(174) <= not(p174_out);
    p174 : perceptron
        Generic map (
            WEIGHTS => "11",
            SHIFT => 6,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p174_in,
            y(0) => p174_out,
            y(1 to 12 - 1) => dummy174
        );


    p175_in <= x(53) & x(130);
    y(175) <= not(p175_out);
    p175 : perceptron
        Generic map (
            WEIGHTS => "01",
            SHIFT => 6,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p175_in,
            y(0) => p175_out,
            y(1 to 12 - 1) => dummy175
        );


    p176_in <= x(49) & x(184) & x(203);
    y(176) <= not(p176_out);
    p176 : perceptron
        Generic map (
            WEIGHTS => "011",
            SHIFT => 6,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p176_in,
            y(0) => p176_out,
            y(1 to 13 - 1) => dummy176
        );


    p177_in <= x(5) & x(166);
    y(177) <= not(p177_out);
    p177 : perceptron
        Generic map (
            WEIGHTS => "00",
            SHIFT => 6,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p177_in,
            y(0) => p177_out,
            y(1 to 12 - 1) => dummy177
        );


    p178_in <= x(80) & x(190);
    y(178) <= not(p178_out);
    p178 : perceptron
        Generic map (
            WEIGHTS => "10",
            SHIFT => 7,
            B => 10,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p178_in,
            y(0) => p178_out,
            y(1 to 13 - 1) => dummy178
        );


    p179_in(0) <= x(226);
    y(179) <= not(p179_out);
    p179 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p179_in,
            y(0) => p179_out,
            y(1 to 12 - 1) => dummy179
        );


    p180_in(0) <= x(80);
    y(180) <= not(p180_out);
    p180 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => 5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p180_in,
            y(0) => p180_out,
            y(1 to 12 - 1) => dummy180
        );


    p181_in <= x(30) & x(33);
    y(181) <= not(p181_out);
    p181 : perceptron
        Generic map (
            WEIGHTS => "10",
            SHIFT => 6,
            B => 9,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p181_in,
            y(0) => p181_out,
            y(1 to 12 - 1) => dummy181
        );


    p182_in <= x(7) & x(40) & x(157);
    y(182) <= not(p182_out);
    p182 : perceptron
        Generic map (
            WEIGHTS => "010",
            SHIFT => 6,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p182_in,
            y(0) => p182_out,
            y(1 to 13 - 1) => dummy182
        );


    p183_in <= x(103) & x(185) & x(253);
    y(183) <= not(p183_out);
    p183 : perceptron
        Generic map (
            WEIGHTS => "001",
            SHIFT => 6,
            B => 5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p183_in,
            y(0) => p183_out,
            y(1 to 13 - 1) => dummy183
        );


    p184_in <= x(107) & x(244);
    y(184) <= not(p184_out);
    p184 : perceptron
        Generic map (
            WEIGHTS => "11",
            SHIFT => 6,
            B => 5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p184_in,
            y(0) => p184_out,
            y(1 to 12 - 1) => dummy184
        );


    p185_in <= x(53) & x(117) & x(195);
    y(185) <= not(p185_out);
    p185 : perceptron
        Generic map (
            WEIGHTS => "101",
            SHIFT => 6,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p185_in,
            y(0) => p185_out,
            y(1 to 13 - 1) => dummy185
        );


    p186_in <= x(58) & x(155);
    y(186) <= not(p186_out);
    p186 : perceptron
        Generic map (
            WEIGHTS => "11",
            SHIFT => 6,
            B => -12,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p186_in,
            y(0) => p186_out,
            y(1 to 12 - 1) => dummy186
        );


    p187_in <= x(32) & x(134);
    y(187) <= not(p187_out);
    p187 : perceptron
        Generic map (
            WEIGHTS => "10",
            SHIFT => 6,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p187_in,
            y(0) => p187_out,
            y(1 to 12 - 1) => dummy187
        );


    p188_in <= x(27) & x(134) & x(166) & x(184) & x(212);
    y(188) <= not(p188_out);
    p188 : perceptron
        Generic map (
            WEIGHTS => "01101",
            SHIFT => 6,
            B => -17,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p188_in,
            y(0) => p188_out,
            y(1 to 14 - 1) => dummy188
        );


    p189_in(0) <= x(105);
    y(189) <= not(p189_out);
    p189 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p189_in,
            y(0) => p189_out,
            y(1 to 12 - 1) => dummy189
        );


    p190_in <= x(29) & x(39);
    y(190) <= not(p190_out);
    p190 : perceptron
        Generic map (
            WEIGHTS => "01",
            SHIFT => 6,
            B => 15,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p190_in,
            y(0) => p190_out,
            y(1 to 12 - 1) => dummy190
        );


    p191_in(0) <= x(190);
    y(191) <= not(p191_out);
    p191 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => -11,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p191_in,
            y(0) => p191_out,
            y(1 to 12 - 1) => dummy191
        );


    p192_in(0) <= x(31);
    y(192) <= not(p192_out);
    p192 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => -10,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p192_in,
            y(0) => p192_out,
            y(1 to 12 - 1) => dummy192
        );


    p193_in(0) <= x(57);
    y(193) <= not(p193_out);
    p193 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p193_in,
            y(0) => p193_out,
            y(1 to 12 - 1) => dummy193
        );


    p194_in(0) <= x(130);
    y(194) <= not(p194_out);
    p194 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p194_in,
            y(0) => p194_out,
            y(1 to 12 - 1) => dummy194
        );


    p195_in(0) <= x(153);
    y(195) <= not(p195_out);
    p195 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => -6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p195_in,
            y(0) => p195_out,
            y(1 to 12 - 1) => dummy195
        );


    p196_in <= x(14) & x(96) & x(250);
    y(196) <= not(p196_out);
    p196 : perceptron
        Generic map (
            WEIGHTS => "001",
            SHIFT => 6,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p196_in,
            y(0) => p196_out,
            y(1 to 13 - 1) => dummy196
        );


    p197_in(0) <= x(73);
    y(197) <= not(p197_out);
    p197 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => -10,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p197_in,
            y(0) => p197_out,
            y(1 to 12 - 1) => dummy197
        );


    p198_in <= x(50) & x(129) & x(235);
    y(198) <= not(p198_out);
    p198 : perceptron
        Generic map (
            WEIGHTS => "001",
            SHIFT => 6,
            B => -6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p198_in,
            y(0) => p198_out,
            y(1 to 13 - 1) => dummy198
        );


    p199_in(0) <= x(9);
    y(199) <= not(p199_out);
    p199 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => 9,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p199_in,
            y(0) => p199_out,
            y(1 to 12 - 1) => dummy199
        );


    p200_in(0) <= x(243);
    y(200) <= not(p200_out);
    p200 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p200_in,
            y(0) => p200_out,
            y(1 to 12 - 1) => dummy200
        );


    p201_in(0) <= x(40);
    y(201) <= not(p201_out);
    p201 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => -7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p201_in,
            y(0) => p201_out,
            y(1 to 12 - 1) => dummy201
        );


    p202_in <= x(32) & x(53);
    y(202) <= not(p202_out);
    p202 : perceptron
        Generic map (
            WEIGHTS => "01",
            SHIFT => 6,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p202_in,
            y(0) => p202_out,
            y(1 to 12 - 1) => dummy202
        );


    p203_in <= x(39) & x(204) & x(235);
    y(203) <= not(p203_out);
    p203 : perceptron
        Generic map (
            WEIGHTS => "101",
            SHIFT => 6,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p203_in,
            y(0) => p203_out,
            y(1 to 13 - 1) => dummy203
        );


    p204_in(0) <= x(177);
    y(204) <= not(p204_out);
    p204 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => 4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p204_in,
            y(0) => p204_out,
            y(1 to 12 - 1) => dummy204
        );


    p205_in <= x(80) & x(235);
    y(205) <= not(p205_out);
    p205 : perceptron
        Generic map (
            WEIGHTS => "01",
            SHIFT => 6,
            B => -8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p205_in,
            y(0) => p205_out,
            y(1 to 12 - 1) => dummy205
        );


    p206_in <= x(19) & x(129) & x(171) & x(177);
    y(206) <= not(p206_out);
    p206 : perceptron
        Generic map (
            WEIGHTS => "1001",
            SHIFT => 6,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p206_in,
            y(0) => p206_out,
            y(1 to 14 - 1) => dummy206
        );


    p207_in <= x(195) & x(228);
    y(207) <= not(p207_out);
    p207 : perceptron
        Generic map (
            WEIGHTS => "10",
            SHIFT => 6,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p207_in,
            y(0) => p207_out,
            y(1 to 12 - 1) => dummy207
        );


    p208_in(0) <= x(32);
    y(208) <= not(p208_out);
    p208 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => 8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p208_in,
            y(0) => p208_out,
            y(1 to 12 - 1) => dummy208
        );


    p209_in <= x(33) & x(38);
    y(209) <= not(p209_out);
    p209 : perceptron
        Generic map (
            WEIGHTS => "01",
            SHIFT => 6,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p209_in,
            y(0) => p209_out,
            y(1 to 12 - 1) => dummy209
        );


    p210_in <= x(177) & x(185) & x(226);
    y(210) <= not(p210_out);
    p210 : perceptron
        Generic map (
            WEIGHTS => "100",
            SHIFT => 6,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p210_in,
            y(0) => p210_out,
            y(1 to 13 - 1) => dummy210
        );


    p211_in <= x(88) & x(110) & x(191);
    y(211) <= not(p211_out);
    p211 : perceptron
        Generic map (
            WEIGHTS => "000",
            SHIFT => 5,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p211_in,
            y(0) => p211_out,
            y(1 to 12 - 1) => dummy211
        );


    p212_in <= x(6) & x(191);
    y(212) <= not(p212_out);
    p212 : perceptron
        Generic map (
            WEIGHTS => "10",
            SHIFT => 6,
            B => -11,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p212_in,
            y(0) => p212_out,
            y(1 to 12 - 1) => dummy212
        );


    p213_in(0) <= x(143);
    y(213) <= not(p213_out);
    p213 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p213_in,
            y(0) => p213_out,
            y(1 to 12 - 1) => dummy213
        );


    p214_in(0) <= x(130);
    y(214) <= not(p214_out);
    p214 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => 4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p214_in,
            y(0) => p214_out,
            y(1 to 12 - 1) => dummy214
        );


    p215_in <= x(165) & x(236);
    y(215) <= not(p215_out);
    p215 : perceptron
        Generic map (
            WEIGHTS => "10",
            SHIFT => 6,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p215_in,
            y(0) => p215_out,
            y(1 to 12 - 1) => dummy215
        );


    p216_in(0) <= x(60);
    y(216) <= not(p216_out);
    p216 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p216_in,
            y(0) => p216_out,
            y(1 to 12 - 1) => dummy216
        );


    p217_in(0) <= x(114);
    y(217) <= not(p217_out);
    p217 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => -6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p217_in,
            y(0) => p217_out,
            y(1 to 12 - 1) => dummy217
        );


    p218_in(0) <= x(164);
    y(218) <= not(p218_out);
    p218 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => -6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p218_in,
            y(0) => p218_out,
            y(1 to 12 - 1) => dummy218
        );


    p219_in(0) <= x(42);
    y(219) <= not(p219_out);
    p219 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => -13,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p219_in,
            y(0) => p219_out,
            y(1 to 12 - 1) => dummy219
        );


    p220_in <= x(117) & x(195) & x(199) & x(249);
    y(220) <= not(p220_out);
    p220 : perceptron
        Generic map (
            WEIGHTS => "0100",
            SHIFT => 6,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p220_in,
            y(0) => p220_out,
            y(1 to 14 - 1) => dummy220
        );


    p221_in <= x(31) & x(195) & x(249);
    y(221) <= not(p221_out);
    p221 : perceptron
        Generic map (
            WEIGHTS => "010",
            SHIFT => 6,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p221_in,
            y(0) => p221_out,
            y(1 to 13 - 1) => dummy221
        );


    p222_in <= x(49) & x(191);
    y(222) <= not(p222_out);
    p222 : perceptron
        Generic map (
            WEIGHTS => "10",
            SHIFT => 6,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p222_in,
            y(0) => p222_out,
            y(1 to 12 - 1) => dummy222
        );


    p223_in <= x(33) & x(65);
    y(223) <= not(p223_out);
    p223 : perceptron
        Generic map (
            WEIGHTS => "11",
            SHIFT => 7,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p223_in,
            y(0) => p223_out,
            y(1 to 13 - 1) => dummy223
        );


    p224_in <= x(144) & x(173) & x(204);
    y(224) <= not(p224_out);
    p224 : perceptron
        Generic map (
            WEIGHTS => "101",
            SHIFT => 6,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p224_in,
            y(0) => p224_out,
            y(1 to 13 - 1) => dummy224
        );


    p225_in <= x(40) & x(68);
    y(225) <= not(p225_out);
    p225 : perceptron
        Generic map (
            WEIGHTS => "11",
            SHIFT => 7,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p225_in,
            y(0) => p225_out,
            y(1 to 13 - 1) => dummy225
        );


    p226_in <= x(80) & x(85) & x(137);
    y(226) <= not(p226_out);
    p226 : perceptron
        Generic map (
            WEIGHTS => "010",
            SHIFT => 6,
            B => -8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p226_in,
            y(0) => p226_out,
            y(1 to 13 - 1) => dummy226
        );


    p227_in <= x(39) & x(239);
    y(227) <= not(p227_out);
    p227 : perceptron
        Generic map (
            WEIGHTS => "01",
            SHIFT => 6,
            B => -12,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p227_in,
            y(0) => p227_out,
            y(1 to 12 - 1) => dummy227
        );


    p228_in <= x(7) & x(88) & x(91) & x(157);
    y(228) <= not(p228_out);
    p228 : perceptron
        Generic map (
            WEIGHTS => "0000",
            SHIFT => 6,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p228_in,
            y(0) => p228_out,
            y(1 to 13 - 1) => dummy228
        );


    p229_in <= x(113) & x(232);
    y(229) <= not(p229_out);
    p229 : perceptron
        Generic map (
            WEIGHTS => "10",
            SHIFT => 6,
            B => 6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p229_in,
            y(0) => p229_out,
            y(1 to 12 - 1) => dummy229
        );


    p230_in(0) <= x(144);
    y(230) <= not(p230_out);
    p230 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => 6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p230_in,
            y(0) => p230_out,
            y(1 to 12 - 1) => dummy230
        );


    p231_in <= x(56) & x(60);
    y(231) <= not(p231_out);
    p231 : perceptron
        Generic map (
            WEIGHTS => "10",
            SHIFT => 6,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p231_in,
            y(0) => p231_out,
            y(1 to 12 - 1) => dummy231
        );


    p232_in <= x(38) & x(177) & x(204) & x(213);
    y(232) <= not(p232_out);
    p232 : perceptron
        Generic map (
            WEIGHTS => "0100",
            SHIFT => 6,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p232_in,
            y(0) => p232_out,
            y(1 to 14 - 1) => dummy232
        );


    p233_in <= x(103) & x(117);
    y(233) <= not(p233_out);
    p233 : perceptron
        Generic map (
            WEIGHTS => "01",
            SHIFT => 7,
            B => 5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p233_in,
            y(0) => p233_out,
            y(1 to 13 - 1) => dummy233
        );


    p234_in(0) <= x(216);
    y(234) <= not(p234_out);
    p234 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => -18,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p234_in,
            y(0) => p234_out,
            y(1 to 12 - 1) => dummy234
        );


    p235_in <= x(33) & x(234);
    y(235) <= not(p235_out);
    p235 : perceptron
        Generic map (
            WEIGHTS => "00",
            SHIFT => 6,
            B => 6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p235_in,
            y(0) => p235_out,
            y(1 to 12 - 1) => dummy235
        );


    p236_in <= x(91) & x(230);
    y(236) <= not(p236_out);
    p236 : perceptron
        Generic map (
            WEIGHTS => "01",
            SHIFT => 6,
            B => 8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p236_in,
            y(0) => p236_out,
            y(1 to 12 - 1) => dummy236
        );


    p237_in <= x(117) & x(121) & x(199);
    y(237) <= not(p237_out);
    p237 : perceptron
        Generic map (
            WEIGHTS => "000",
            SHIFT => 6,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p237_in,
            y(0) => p237_out,
            y(1 to 13 - 1) => dummy237
        );


    p238_in <= x(39) & x(66) & x(133);
    y(238) <= not(p238_out);
    p238 : perceptron
        Generic map (
            WEIGHTS => "010",
            SHIFT => 5,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p238_in,
            y(0) => p238_out,
            y(1 to 12 - 1) => dummy238
        );


    p239_in <= x(6) & x(53) & x(140);
    y(239) <= not(p239_out);
    p239 : perceptron
        Generic map (
            WEIGHTS => "001",
            SHIFT => 6,
            B => 5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p239_in,
            y(0) => p239_out,
            y(1 to 13 - 1) => dummy239
        );


    p240_in <= x(31) & x(126);
    y(240) <= not(p240_out);
    p240 : perceptron
        Generic map (
            WEIGHTS => "10",
            SHIFT => 6,
            B => 7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p240_in,
            y(0) => p240_out,
            y(1 to 12 - 1) => dummy240
        );


    p241_in(0) <= x(201);
    y(241) <= not(p241_out);
    p241 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => 7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p241_in,
            y(0) => p241_out,
            y(1 to 12 - 1) => dummy241
        );


    p242_in <= x(45) & x(100) & x(185) & x(242);
    y(242) <= not(p242_out);
    p242 : perceptron
        Generic map (
            WEIGHTS => "1100",
            SHIFT => 6,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p242_in,
            y(0) => p242_out,
            y(1 to 14 - 1) => dummy242
        );


    p243_in(0) <= x(60);
    y(243) <= not(p243_out);
    p243 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => -6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p243_in,
            y(0) => p243_out,
            y(1 to 12 - 1) => dummy243
        );


    p244_in <= x(9) & x(126) & x(141) & x(195);
    y(244) <= not(p244_out);
    p244 : perceptron
        Generic map (
            WEIGHTS => "0111",
            SHIFT => 6,
            B => -15,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p244_in,
            y(0) => p244_out,
            y(1 to 13 - 1) => dummy244
        );


    p245_in <= x(65) & x(174);
    y(245) <= not(p245_out);
    p245 : perceptron
        Generic map (
            WEIGHTS => "01",
            SHIFT => 6,
            B => -8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p245_in,
            y(0) => p245_out,
            y(1 to 12 - 1) => dummy245
        );


    p246_in <= x(32) & x(53) & x(132) & x(140) & x(184) & x(189);
    y(246) <= not(p246_out);
    p246 : perceptron
        Generic map (
            WEIGHTS => "000101",
            SHIFT => 5,
            B => 4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p246_in,
            y(0) => p246_out,
            y(1 to 13 - 1) => dummy246
        );


    p247_in(0) <= x(216);
    y(247) <= not(p247_out);
    p247 : perceptron
        Generic map (
            WEIGHTS => "1",
            SHIFT => 7,
            B => -18,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p247_in,
            y(0) => p247_out,
            y(1 to 12 - 1) => dummy247
        );


    p248_in <= x(96) & x(143);
    y(248) <= not(p248_out);
    p248 : perceptron
        Generic map (
            WEIGHTS => "00",
            SHIFT => 6,
            B => -12,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p248_in,
            y(0) => p248_out,
            y(1 to 12 - 1) => dummy248
        );


    p249_in(0) <= x(177);
    y(249) <= not(p249_out);
    p249 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => -6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p249_in,
            y(0) => p249_out,
            y(1 to 12 - 1) => dummy249
        );


    p250_in <= x(132) & x(177) & x(189) & x(201) & x(251) & x(252);
    y(250) <= not(p250_out);
    p250 : perceptron
        Generic map (
            WEIGHTS => "010000",
            SHIFT => 6,
            B => 9,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p250_in,
            y(0) => p250_out,
            y(1 to 14 - 1) => dummy250
        );


    p251_in(0) <= x(94);
    y(251) <= not(p251_out);
    p251 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p251_in,
            y(0) => p251_out,
            y(1 to 12 - 1) => dummy251
        );


    p252_in <= x(0) & x(32) & x(236) & x(251);
    y(252) <= not(p252_out);
    p252 : perceptron
        Generic map (
            WEIGHTS => "0101",
            SHIFT => 6,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p252_in,
            y(0) => p252_out,
            y(1 to 13 - 1) => dummy252
        );


    p253_in(0) <= x(100);
    y(253) <= not(p253_out);
    p253 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => 11,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p253_in,
            y(0) => p253_out,
            y(1 to 12 - 1) => dummy253
        );


    p254_in(0) <= x(46);
    y(254) <= not(p254_out);
    p254 : perceptron
        Generic map (
            WEIGHTS => "0",
            SHIFT => 7,
            B => 5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p254_in,
            y(0) => p254_out,
            y(1 to 12 - 1) => dummy254
        );


    p255_in <= x(6) & x(78);
    y(255) <= not(p255_out);
    p255 : perceptron
        Generic map (
            WEIGHTS => "10",
            SHIFT => 7,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p255_in,
            y(0) => p255_out,
            y(1 to 13 - 1) => dummy255
        );



end layer_4;

architecture layer_5 of layer is

    Component perceptron
    Generic (
        WEIGHTS : STD_LOGIC_VECTOR := (others => '0');
        SHIFT : Integer;     -- number of shift (left + or right -)
        B : Integer;          -- bias of batch norm
        BATCH_POSITIVE : Boolean    
    );
    Port ( 
        x : in STD_LOGIC_VECTOR;
        y : out STD_LOGIC_VECTOR
   );
    end component;
    
    -- Signals
    signal p0_in : STD_LOGIC_VECTOR(0 to 95 - 1);
	signal p0_out : STD_LOGIC;
	signal p1_in : STD_LOGIC_VECTOR(0 to 105 - 1);
	signal p1_out : STD_LOGIC;
	signal p2_in : STD_LOGIC_VECTOR(0 to 100 - 1);
	signal p2_out : STD_LOGIC;
	signal p3_in : STD_LOGIC_VECTOR(0 to 79 - 1);
	signal p3_out : STD_LOGIC;
	signal p4_in : STD_LOGIC_VECTOR(0 to 89 - 1);
	signal p4_out : STD_LOGIC;
	signal p5_in : STD_LOGIC_VECTOR(0 to 86 - 1);
	signal p5_out : STD_LOGIC;
	signal p6_in : STD_LOGIC_VECTOR(0 to 103 - 1);
	signal p6_out : STD_LOGIC;
	signal p7_in : STD_LOGIC_VECTOR(0 to 100 - 1);
	signal p7_out : STD_LOGIC;
	signal p8_in : STD_LOGIC_VECTOR(0 to 66 - 1);
	signal p8_out : STD_LOGIC;
	signal p9_in : STD_LOGIC_VECTOR(0 to 83 - 1);
	signal p9_out : STD_LOGIC;
	
    
    -- Dummies
     

begin

    
    p0_in <= x(3) & x(4) & x(5) & x(6) & x(7) & x(17) & x(21) & x(29) & x(32) & x(35) & x(38) & x(39) & x(40) & x(47) & x(53) & x(54) & x(59) & x(66) & x(67) & x(72) & x(73) & x(74) & x(76) & x(79) & x(81) & x(87) & x(88) & x(92) & x(95) & x(96) & x(99) & x(100) & x(101) & x(104) & x(105) & x(106) & x(111) & x(113) & x(114) & x(115) & x(122) & x(126) & x(129) & x(130) & x(132) & x(133) & x(134) & x(135) & x(136) & x(140) & x(143) & x(144) & x(146) & x(147) & x(148) & x(150) & x(155) & x(156) & x(163) & x(164) & x(165) & x(167) & x(171) & x(172) & x(173) & x(174) & x(175) & x(178) & x(180) & x(184) & x(186) & x(189) & x(191) & x(192) & x(193) & x(195) & x(200) & x(202) & x(205) & x(211) & x(212) & x(213) & x(214) & x(217) & x(218) & x(221) & x(223) & x(228) & x(235) & x(236) & x(237) & x(239) & x(243) & x(246) & x(254);
    p0 : perceptron
        Generic map (
            WEIGHTS => "00001000111110111000110010111010111001111001100110010011011101001111111011111000011011000011011",
            SHIFT => -3,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p0_in,
            y => y(0 to 8)
        );


    p1_in <= x(2) & x(3) & x(6) & x(8) & x(9) & x(10) & x(13) & x(14) & x(15) & x(19) & x(20) & x(21) & x(22) & x(28) & x(30) & x(31) & x(36) & x(40) & x(42) & x(44) & x(45) & x(48) & x(50) & x(51) & x(52) & x(54) & x(56) & x(59) & x(60) & x(65) & x(67) & x(69) & x(71) & x(72) & x(77) & x(79) & x(80) & x(81) & x(82) & x(86) & x(88) & x(89) & x(91) & x(92) & x(102) & x(106) & x(107) & x(110) & x(111) & x(113) & x(119) & x(120) & x(121) & x(123) & x(124) & x(128) & x(129) & x(130) & x(132) & x(134) & x(137) & x(145) & x(149) & x(150) & x(154) & x(155) & x(158) & x(159) & x(160) & x(165) & x(166) & x(168) & x(169) & x(171) & x(172) & x(175) & x(179) & x(184) & x(185) & x(190) & x(191) & x(192) & x(193) & x(194) & x(195) & x(197) & x(207) & x(209) & x(212) & x(214) & x(217) & x(218) & x(219) & x(220) & x(221) & x(224) & x(225) & x(227) & x(229) & x(235) & x(237) & x(238) & x(248) & x(249) & x(251);
    p1 : perceptron
        Generic map (
            WEIGHTS => "011011101101000110010010001010110101000001001101101011011001111001010101011000000001000100100001010101000",
            SHIFT => -3,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p1_in,
            y => y(9 to 17)
        );


    p2_in <= x(0) & x(3) & x(4) & x(7) & x(8) & x(10) & x(13) & x(17) & x(19) & x(22) & x(25) & x(26) & x(27) & x(28) & x(31) & x(35) & x(38) & x(39) & x(40) & x(41) & x(42) & x(47) & x(50) & x(53) & x(54) & x(55) & x(57) & x(58) & x(61) & x(63) & x(68) & x(71) & x(74) & x(76) & x(78) & x(79) & x(81) & x(82) & x(83) & x(89) & x(93) & x(99) & x(100) & x(102) & x(107) & x(112) & x(113) & x(116) & x(121) & x(123) & x(126) & x(133) & x(134) & x(136) & x(138) & x(143) & x(144) & x(145) & x(146) & x(149) & x(152) & x(157) & x(163) & x(164) & x(165) & x(167) & x(168) & x(170) & x(171) & x(174) & x(177) & x(180) & x(185) & x(193) & x(195) & x(202) & x(203) & x(204) & x(205) & x(206) & x(207) & x(208) & x(209) & x(219) & x(220) & x(221) & x(223) & x(224) & x(231) & x(233) & x(235) & x(236) & x(238) & x(242) & x(244) & x(248) & x(251) & x(252) & x(253) & x(254);
    p2 : perceptron
        Generic map (
            WEIGHTS => "0001100010001111010100011100011001100101100101101100111101011000011110010110000100110001011111001111",
            SHIFT => -3,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p2_in,
            y => y(18 to 26)
        );


    p3_in <= x(11) & x(17) & x(19) & x(20) & x(22) & x(23) & x(24) & x(25) & x(26) & x(31) & x(33) & x(37) & x(42) & x(47) & x(48) & x(51) & x(54) & x(57) & x(59) & x(61) & x(62) & x(64) & x(78) & x(79) & x(80) & x(82) & x(83) & x(86) & x(93) & x(96) & x(105) & x(113) & x(114) & x(115) & x(118) & x(123) & x(124) & x(125) & x(126) & x(130) & x(132) & x(133) & x(149) & x(156) & x(158) & x(165) & x(166) & x(167) & x(168) & x(171) & x(177) & x(178) & x(180) & x(182) & x(184) & x(187) & x(188) & x(189) & x(196) & x(198) & x(199) & x(201) & x(202) & x(203) & x(205) & x(217) & x(218) & x(228) & x(229) & x(230) & x(233) & x(234) & x(237) & x(238) & x(244) & x(247) & x(248) & x(254) & x(255);
    p3 : perceptron
        Generic map (
            WEIGHTS => "0000010111110101011001100000001010110011101100111101001011001110010011001100011",
            SHIFT => -3,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p3_in,
            y => y(27 to 35)
        );


    p4_in <= x(22) & x(28) & x(30) & x(31) & x(32) & x(35) & x(41) & x(42) & x(43) & x(44) & x(49) & x(53) & x(55) & x(63) & x(71) & x(73) & x(76) & x(79) & x(80) & x(86) & x(87) & x(89) & x(97) & x(101) & x(103) & x(105) & x(106) & x(107) & x(108) & x(109) & x(110) & x(112) & x(114) & x(116) & x(122) & x(123) & x(125) & x(128) & x(130) & x(133) & x(134) & x(137) & x(139) & x(140) & x(144) & x(145) & x(147) & x(149) & x(150) & x(151) & x(152) & x(154) & x(156) & x(157) & x(158) & x(161) & x(162) & x(164) & x(168) & x(170) & x(173) & x(174) & x(176) & x(178) & x(179) & x(183) & x(190) & x(191) & x(192) & x(195) & x(203) & x(205) & x(209) & x(210) & x(214) & x(220) & x(222) & x(224) & x(226) & x(227) & x(228) & x(230) & x(231) & x(237) & x(238) & x(242) & x(248) & x(249) & x(251);
    p4 : perceptron
        Generic map (
            WEIGHTS => "11000001110001101111100100111101010010010111001001010111100000100011111100010010101000110",
            SHIFT => -3,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p4_in,
            y => y(36 to 44)
        );


    p5_in <= x(0) & x(1) & x(12) & x(13) & x(14) & x(15) & x(17) & x(20) & x(24) & x(26) & x(28) & x(33) & x(34) & x(37) & x(39) & x(48) & x(52) & x(59) & x(62) & x(64) & x(65) & x(70) & x(73) & x(74) & x(87) & x(94) & x(95) & x(98) & x(99) & x(104) & x(111) & x(113) & x(114) & x(115) & x(116) & x(120) & x(122) & x(125) & x(127) & x(130) & x(134) & x(135) & x(140) & x(148) & x(151) & x(152) & x(153) & x(154) & x(156) & x(158) & x(159) & x(160) & x(162) & x(166) & x(173) & x(174) & x(177) & x(181) & x(182) & x(185) & x(186) & x(191) & x(194) & x(198) & x(199) & x(201) & x(203) & x(210) & x(214) & x(217) & x(219) & x(220) & x(221) & x(223) & x(226) & x(227) & x(228) & x(233) & x(234) & x(236) & x(237) & x(241) & x(244) & x(247) & x(253) & x(254);
    p5 : perceptron
        Generic map (
            WEIGHTS => "10110110011111000101001101111100111110010101100110011101100111110111110111000000101000",
            SHIFT => -3,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p5_in,
            y => y(45 to 53)
        );


    p6_in <= x(0) & x(1) & x(5) & x(7) & x(8) & x(9) & x(10) & x(15) & x(19) & x(21) & x(26) & x(27) & x(28) & x(33) & x(34) & x(38) & x(42) & x(53) & x(55) & x(56) & x(58) & x(61) & x(67) & x(69) & x(71) & x(73) & x(79) & x(80) & x(82) & x(86) & x(87) & x(88) & x(90) & x(93) & x(94) & x(99) & x(102) & x(106) & x(107) & x(111) & x(112) & x(116) & x(120) & x(121) & x(122) & x(123) & x(124) & x(125) & x(126) & x(127) & x(131) & x(132) & x(134) & x(142) & x(144) & x(145) & x(146) & x(148) & x(149) & x(150) & x(154) & x(155) & x(156) & x(159) & x(160) & x(164) & x(170) & x(174) & x(176) & x(180) & x(182) & x(185) & x(191) & x(193) & x(194) & x(195) & x(196) & x(197) & x(198) & x(206) & x(207) & x(208) & x(209) & x(215) & x(218) & x(219) & x(220) & x(221) & x(222) & x(226) & x(230) & x(233) & x(235) & x(237) & x(241) & x(244) & x(245) & x(248) & x(249) & x(250) & x(252) & x(253) & x(255);
    p6 : perceptron
        Generic map (
            WEIGHTS => "0011100110011001011001111111110101000110001000110000010011001001011001101111111101000100101100100111010",
            SHIFT => -3,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p6_in,
            y => y(54 to 62)
        );


    p7_in <= x(3) & x(4) & x(6) & x(8) & x(12) & x(14) & x(18) & x(20) & x(21) & x(22) & x(24) & x(27) & x(28) & x(32) & x(35) & x(41) & x(42) & x(43) & x(44) & x(46) & x(47) & x(48) & x(49) & x(52) & x(55) & x(58) & x(60) & x(63) & x(65) & x(67) & x(68) & x(69) & x(71) & x(73) & x(74) & x(76) & x(81) & x(85) & x(88) & x(93) & x(99) & x(103) & x(108) & x(113) & x(114) & x(119) & x(120) & x(121) & x(124) & x(125) & x(126) & x(129) & x(133) & x(135) & x(136) & x(137) & x(140) & x(141) & x(142) & x(144) & x(150) & x(151) & x(152) & x(155) & x(156) & x(157) & x(158) & x(159) & x(162) & x(168) & x(170) & x(173) & x(174) & x(179) & x(180) & x(183) & x(184) & x(185) & x(187) & x(188) & x(194) & x(198) & x(200) & x(201) & x(204) & x(205) & x(208) & x(211) & x(212) & x(216) & x(217) & x(218) & x(223) & x(225) & x(226) & x(230) & x(231) & x(236) & x(243) & x(245);
    p7 : perceptron
        Generic map (
            WEIGHTS => "0010010111100100100101010110100010101100100101010110101000011001011000011000011000001100010101101011",
            SHIFT => -3,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p7_in,
            y => y(63 to 71)
        );


    p8_in <= x(1) & x(3) & x(16) & x(17) & x(23) & x(25) & x(27) & x(35) & x(36) & x(37) & x(38) & x(41) & x(47) & x(51) & x(52) & x(55) & x(58) & x(61) & x(62) & x(66) & x(68) & x(69) & x(75) & x(81) & x(83) & x(84) & x(87) & x(89) & x(95) & x(98) & x(100) & x(101) & x(102) & x(104) & x(105) & x(114) & x(122) & x(125) & x(137) & x(140) & x(148) & x(154) & x(156) & x(157) & x(168) & x(171) & x(172) & x(175) & x(180) & x(184) & x(186) & x(187) & x(188) & x(196) & x(205) & x(209) & x(213) & x(226) & x(230) & x(234) & x(236) & x(237) & x(247) & x(248) & x(252) & x(254);
    p8 : perceptron
        Generic map (
            WEIGHTS => "110100010001110101111010101101100111100100101001111011010001111100",
            SHIFT => -2,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p8_in,
            y => y(72 to 81)
        );


    p9_in <= x(1) & x(7) & x(12) & x(19) & x(22) & x(27) & x(28) & x(30) & x(31) & x(32) & x(35) & x(41) & x(42) & x(43) & x(44) & x(53) & x(55) & x(58) & x(63) & x(64) & x(66) & x(67) & x(71) & x(73) & x(79) & x(80) & x(86) & x(87) & x(91) & x(95) & x(97) & x(101) & x(102) & x(104) & x(105) & x(106) & x(110) & x(120) & x(125) & x(127) & x(129) & x(130) & x(131) & x(133) & x(135) & x(139) & x(140) & x(141) & x(145) & x(147) & x(148) & x(149) & x(150) & x(151) & x(156) & x(158) & x(161) & x(165) & x(170) & x(171) & x(178) & x(179) & x(192) & x(194) & x(203) & x(205) & x(209) & x(210) & x(211) & x(213) & x(216) & x(218) & x(221) & x(224) & x(226) & x(228) & x(229) & x(231) & x(232) & x(238) & x(242) & x(248) & x(249);
    p9 : perceptron
        Generic map (
            WEIGHTS => "10001001000010000100111011111010000000111011001100001001110001101101100110111010110",
            SHIFT => -3,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p9_in,
            y => y(82 to 90)
        );



end layer_5;
